*simulator lang=spice


*** .LIB MOS ***
.SUBCKT NENHHP_S D G S B l=0 wpf=0 as=0 ad=0 ps=0 pd=0 nrs=0 nrd=0 simM=1 sa=0 sb=0 sc=0 sca=0 scb=0 scc=0 mcm_NENHHP_vth0=0 mcm_NENHHP_u0=0
** Pelgrom Scaling parameter **
.param mcmScale='1/sqrt(l*wpf)*1/sqrt(simM)'

.flat M0
M0 D G S B NENHHP  l=l w=wpf as=as ad=ad ps=ps pd=pd nrs=nrs nrd=nrd
+ m=simM sa=sa sb=sb sc=sc sca=sca scb=scb scc=scc

.MODEL NENHHP.001 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.362+dvth0n001_hp+(mcm_NENHHP_vth0*mcmScale)'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.13
+NFACTOR = 2.25
+ETA0 = 0.12
+ETAB = -0.1
+U0 = '(0.024*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '115000*dvsatfactorn_hp'
+A0 = 1
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0101
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1977
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+LVTH0 = '0.0+dlvth0n001_hp'
+WVTH0 = '0.0+dwvth0n001_hp'
+PVTH0 = '0.0+dpvth0n001_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.101 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.35948434+dvth0n101_hp+(mcm_NENHHP_vth0*mcmScale)'
+WVTH0 = '2.4975463e-08+dwvth0n101_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1347689*dk2factorn_hp'
+WK2 = '-5.1934405e-08*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.11828233
+WVOFF = -1.1633307e-07
+NFACTOR = 2.25
+ETA0 = 0.10744535
+WETA0 = 1.2464257e-07
+ETAB = -0.1
+U0 = '(0.022326047*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+WU0 = '1.661901e-08*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '110815.12*dvsatfactorn_hp'
+WVSAT = '0.041547524*dvsatfactorn_hp'
+A0 = 1
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.012554651
+WKETA = 1.2464257e-07
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010120924
+WAIGC = -2.0773762e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.19686302
+WKT1 = -8.3095048e-09
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4237545
+WUTE = -3.6977296e-07
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+LVTH0 = '0.0+dlvth0n101_hp'
+PVTH0 = '0.0+dpvth0n101_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.201 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.36855982+dvth0n201_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.1631657e-10+dlvth0n201_hp'
+WVTH0 = '-1.6066231e-09+dwvth0n201_hp'
+PVTH0 = '1.8051912e-15+dpvth0n201_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.15640403*dk2factorn_hp'
+LK2 = '2.4230944e-10*dk2factorn_hp'
+WK2 = '1.1434914e-08*dk2factorn_hp'
+PK2 = '-7.0972435e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.17938279
+LVOFF = 1.3483854e-09
+WVOFF = 6.2630202e-08
+PVOFF = -3.9494209e-15
+NFACTOR = 2.25
+ETA0 = 0.17584233
+LETA0 = -1.23578e-09
+WETA0 = -7.5692173e-08
+PETA0 = 3.6195997e-15
+ETAB = -0.1
+U0 = '(0.028819034*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.3615699e-11*du0factorn_hp'
+WU0 = '-2.3989511e-09*du0factorn_hp'
+PU0 = '1.2775038e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '129560.44*dvsatfactorn_hp'
+LVSAT = '-0.00021808038*dvsatfactorn_hp'
+WVSAT = '-0.013357537*dvsatfactorn_hp'
+PVSAT = '6.3875743e-10*dvsatfactorn_hp'
+A0 = 0.73834768
+LA0 = 1.6961698e-08
+WA0 = 7.6637963e-07
+PA0 = -4.9680815e-14
+AGS = 1.1013425
+LAGS = -4.8462001e-09
+WAGS = -2.9683229e-07
+PAGS = 1.419452e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.024932877
+LKETA = 2.4230982e-10
+WKETA = 1.4841603e-08
+PKETA = -7.0972545e-16
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010020516
+LAIGC = 3.6346604e-12
+WAIGC = 8.6358218e-11
+PAIGC = -1.064592e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5971712
+LUTE = 3.3680993e-09
+WUTE = 1.3816453e-07
+PUTE = -9.8651629e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.301 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.25319942+dvth0n301_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '7.650598e-09+dlvth0n301_hp'
+WVTH0 = '1.0567855e-07+dwvth0n301_hp'
+PVTH0 = '-5.8830393e-15+dpvth0n301_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.2143025*dk2factorn_hp'
+LK2 = '3.2506696e-09*dk2factorn_hp'
+WK2 = '6.5280487e-08*dk2factorn_hp'
+PK2 = '-3.5074993e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0032938639
+LCDSCB = -3.8393739e-10
+WCDSCB = -5.8532935e-09
+PCDSCB = 3.5706178e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.11259084
+LVOFF = -2.8408078e-09
+WVOFF = 5.1368066e-10
+PVOFF = -5.3471185e-17
+NFACTOR = 4.0564813
+LNFACTOR = -8.6385934e-08
+WNFACTOR = -1.6800276e-06
+PNFACTOR = 8.0338919e-14
+ETA0 = 0.28922131
+LETA0 = -4.5419602e-09
+WETA0 = -1.8113463e-07
+PETA0 = 6.6943472e-15
+ETAB = -0.1
+U0 = '(0.04144366*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.0798016e-10*du0factorn_hp'
+WU0 = '-1.4139853e-08*du0factorn_hp'
+PU0 = '7.4560933e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 1.5383651e-27
+LUC = -8.4022855e-35
+WUC = -1.6340706e-33
+PUC = 7.8141255e-41
+EU = 2.9
+VSAT = '109841.02*dvsatfactorn_hp'
+LVSAT = '0.00068342004*dvsatfactorn_hp'
+WVSAT = '0.0049815265*dvsatfactorn_hp'
+PVSAT = '-1.9963795e-10*dvsatfactorn_hp'
+A0 = 1.2797015
+LA0 = -1.0494602e-08
+WA0 = 2.6292059e-07
+PA0 = -2.4146455e-14
+AGS = 0.59320536
+LAGS = 1.945292e-08
+WAGS = 1.7573528e-07
+PAGS = -8.4036613e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.050339716
+LKETA = -9.7264523e-10
+WKETA = -8.7867574e-09
+PKETA = 4.2018274e-16
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0093013289
+LAIGC = 3.7241815e-11
+WAIGC = 7.5520239e-10
+PAIGC = -4.1900574e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.20772887
+LKT1 = 3.8394077e-10
+WKT1 = 7.466853e-09
+PKT1 = -3.5706491e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -2.189973
+LUTE = 3.2360749e-08
+WUTE = 6.8947017e-07
+PUTE = -3.6828327e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.401 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.59478745+dvth0n401_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.044021e-08+dlvth0n401_hp'
+WVTH0 = '-4.1887478e-08+dwvth0n401_hp'
+PVTH0 = '1.9321898e-15+dpvth0n401_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '0.0073189607*dk2factorn_hp'
+LK2 = '-8.2402927e-09*dk2factorn_hp'
+WK2 = '-3.0459984e-08*dk2factorn_hp'
+PK2 = '1.4565964e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.015705601
+LCDSCB = 7.367335e-10
+WCDSCB = 2.3544754e-09
+PCDSCB = -1.2706805e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.080273192
+LVOFF = -4.709774e-09
+WVOFF = -1.3447541e-08
+PVOFF = 7.5392222e-16
+NFACTOR = -1.0161072
+LNFACTOR = 1.6456316e-07
+WNFACTOR = 5.1133064e-07
+PNFACTOR = -2.807109e-14
+ETA0 = -0.25975293
+LETA0 = 1.846252e-08
+WETA0 = 5.6022245e-08
+PETA0 = -3.2435881e-15
+ETAB = -0.1
+U0 = '(-0.0058703526*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.7153203e-09*du0factorn_hp'
+WU0 = '6.2998003e-09*du0factorn_hp'
+PU0 = '-3.0125645e-16*du0factorn_hp'
+UA = -5.0772913e-28
+WUA = 3.1109579e-34
+UB = 1e-19
+UC = -3.5023591e-27
+LUC = 1.5702458e-34
+WUC = 5.4352228e-34
+PUC = -2.5991235e-41
+EU = 2.9
+VSAT = '109262.62*dvsatfactorn_hp'
+LVSAT = '0.00026419528*dvsatfactorn_hp'
+WVSAT = '0.0052313971*dvsatfactorn_hp'
+PVSAT = '-1.8532859e-11*dvsatfactorn_hp'
+A0 = 3.0013844
+LA0 = -1.1291387e-07
+WA0 = -4.8084642e-07
+PA0 = 2.0098669e-14
+AGS = 0.7013625
+LAGS = -1.9230808e-08
+WAGS = 1.290114e-07
+PAGS = 8.3077092e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03274048
+LKETA = -8.0128283e-10
+WKETA = -1.1838874e-09
+PKETA = 3.4615418e-16
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.011659719
+LAIGC = -1.0066082e-10
+WAIGC = -2.6362195e-10
+PAIGC = 1.7673363e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.18395835
+LKT1 = -7.5276575e-10
+WKT1 = -2.8020139e-09
+PKT1 = 1.339923e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = 0.064448897
+LUTE = -8.7727112e-08
+WUTE = -2.8444009e-07
+PUTE = 1.5049629e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.501 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.38729287+dvth0n501_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '7.3363057e-10+dlvth0n501_hp'
+WVTH0 = '-4.9534428e-09+dwvth0n501_hp'
+PVTH0 = '-5.6753861e-17+dpvth0n501_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.15671336*dk2factorn_hp'
+LK2 = '-1.2259846e-10*dk2factorn_hp'
+WK2 = '-1.2622308e-09*dk2factorn_hp'
+PK2 = '1.1646853e-17*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0032763619
+LCDSCB = 6.1035625e-11
+WCDSCB = 1.4207083e-10
+PCDSCB = -6.7938273e-18
+CDSCD = 0
+CIT = 0
+VOFF = -0.1651638
+LVOFF = -5.7691437e-10
+WVOFF = 1.6629871e-09
+PVOFF = 1.8273198e-17
+NFACTOR = 1.9463275
+LNFACTOR = 1.3513364e-08
+WNFACTOR = -1.5982746e-08
+PNFACTOR = -1.184226e-15
+ETA0 = 0.014894253
+LETA0 = 5.1494479e-10
+WETA0 = 7.135046e-09
+PETA0 = -4.8919755e-17
+ETAB = -0.1
+U0 = '(0.023753134*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.5056466e-11*du0factorn_hp'
+WU0 = '1.0268197e-09*du0factorn_hp'
+PU0 = '-3.8949375e-19*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -6.1924858e-28
+LUC = 2.3604086e-35
+WUC = 3.0328615e-35
+PUC = -2.2423882e-42
+EU = 2.9
+VSAT = '111003.68*dvsatfactorn_hp'
+LVSAT = '0.00022336804*dvsatfactorn_hp'
+WVSAT = '0.0049214873*dvsatfactorn_hp'
+PVSAT = '-1.1265612e-11*dvsatfactorn_hp'
+A0 = 0.3
+AGS = 1.0702848
+LAGS = 4.445898e-08
+WAGS = 6.3343227e-08
+PAGS = -3.0290731e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.11317974
+LKETA = 2.4521185e-09
+WKETA = -1.5502075e-08
+PKETA = -2.3295126e-16
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010315199
+LAIGC = -7.8442181e-13
+WAIGC = -2.4297437e-11
+PAIGC = -1.0463519e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.2002016
+LKT1 = 2.3986392e-11
+WKT1 = 8.9284352e-11
+PKT1 = -4.2695777e-18
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4699889
+LUTE = -6.2171294e-09
+WUTE = -1.1310157e-08
+PUTE = 5.4085168e-16
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.601 NMOS
+LMIN = '9.00000000e-08+lminoffsetn_hp'
+LMAX = '9.30000000e-08+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.6333514+dvth0n601_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.3722016e-08+dlvth0n601_hp'
+WVTH0 = '-2.8329003e-08+dwvth0n601_hp'
+PVTH0 = '1.3165326e-15+dpvth0n601_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.198*dk2factorn_hp'
+WK2 = '2.66e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0039673417
+LCDSCB = -3.9817718e-11
+WCDSCB = 2.0771392e-10
+PCDSCB = 2.7872403e-18
+CDSCD = 0
+CIT = 0
+VOFF = -0.33873734
+LVOFF = 6.6505695e-09
+WVOFF = 1.8152474e-08
+PVOFF = -6.6833777e-16
+NFACTOR = 4.551601
+LNFACTOR = -1.9183476e-07
+WNFACTOR = -2.6348373e-07
+PNFACTOR = 1.8323846e-14
+ETA0 = 0.74053748
+LETA0 = -3.2447662e-08
+WETA0 = -6.1801061e-08
+PETA0 = 3.0825279e-15
+ETAB = -0.1
+U0 = '(0.0054163917*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.2595985e-10*du0factorn_hp'
+WU0 = '2.7688102e-09*du0factorn_hp'
+PU0 = '3.2957057e-17*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -3e-28
+EU = 2.9
+VSAT = '186307.86*dvsatfactorn_hp'
+LVSAT = '-0.007713742*dvsatfactorn_hp'
+WVSAT = '-0.00223241*dvsatfactorn_hp'
+PVSAT = '7.4275985e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = 1.0008114
+LAGS = 4.77812e-08
+WAGS = 6.9943203e-08
+PAGS = -3.344684e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.20445157
+LKETA = -1.2167874e-08
+WKETA = -2.4172899e-08
+PKETA = 1.155948e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0099162412
+LAIGC = 9.4486658e-13
+WAIGC = 1.3603538e-11
+PAIGC = -2.6891758e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1980347
+LKT1 = -7.963482e-11
+WKT1 = -1.1657125e-10
+PKT1 = 5.5744374e-18
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -2.694708
+LUTE = 7.9128137e-08
+WUTE = 1.0503816e-07
+PUTE = -7.5669486e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = -42931.162
+LAT = 0.0026363722
+WAT = 0.0088284604
+PAT = -2.5045536e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.002 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.48815265+dvth0n002_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.4110775e-09+dlvth0n002_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0040084851
+LCDSCB = -3.5617121e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.038889726
+LVOFF = -4.6302241e-09
+NFACTOR = 2.25
+ETA0 = -0.027178176
+LETA0 = 7.4795949e-09
+ETAB = -0.1
+U0 = '(0.02960679*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.8493708e-10*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '79957.627*dvsatfactorn_hp'
+LVSAT = '0.0017808534*dvsatfactorn_hp'
+A0 = 4.5042425
+LA0 = -1.7808561e-07
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.21025454
+LKETA = -1.0685136e-08
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.00988975
+LAIGC = 1.0684906e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21171684
+LKT1 = 7.1233598e-10
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n002_hp'
+PVTH0 = '0.0+dpvth0n002_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.102 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.5384304+dvth0n102_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-9.0940388e-09+dlvth0n102_hp'
+WVTH0 = '-4.9915755e-07+dwvth0n102_hp'
+PVTH0 = '2.663644e-14+dpvth0n102_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1347689*dk2factorn_hp'
+WK2 = '-5.1934405e-08*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0069414545
+LCDSCB = -5.0522472e-10
+WCDSCB = -2.911852e-08
+PCDSCB = 1.4798032e-15
+CDSCD = 0
+CIT = 0
+VOFF = 0.010956537
+LVOFF = -6.567919e-09
+WVOFF = -4.948737e-07
+PVOFF = 1.9237435e-14
+NFACTOR = 2.25
+ETA0 = -0.10132518
+LETA0 = 1.0609718e-08
+WETA0 = 7.3613145e-07
+PETA0 = -3.1075865e-14
+ETAB = -0.1
+U0 = '(0.030279213*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.0417993e-10*du0factorn_hp'
+WU0 = '-6.6758153e-09*du0factorn_hp'
+PU0 = '1.183843e-15*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '61107.919*dvsatfactorn_hp'
+LVSAT = '0.0025261198*dvsatfactorn_hp'
+WVSAT = '0.18713991*dvsatfactorn_hp'
+PVSAT = '-7.3990048e-09*dvsatfactorn_hp'
+A0 = 5.9707272
+LA0 = -2.5261236e-07
+WA0 = -1.455926e-05
+PA0 = 7.399016e-13
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.28568897
+LKETA = -1.5156741e-08
+WKETA = -7.48913e-07
+PKETA = 4.4394094e-14
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0098226872
+LAIGC = 1.5156414e-11
+WAIGC = 6.6579911e-10
+PAIGC = -4.4393137e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21674575
+LKT1 = 1.0104403e-09
+WKT1 = 4.9927009e-08
+PKT1 = -2.9595796e-15
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4237545
+WUTE = -3.6977296e-07
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.202 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.43002708+dvth0n202_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-3.7400825e-09+dlvth0n202_hp'
+WVTH0 = '-1.8164422e-07+dwvth0n202_hp'
+PVTH0 = '1.0954702e-14+dpvth0n202_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.18057033*dk2factorn_hp'
+LK2 = '1.4704408e-09*dk2factorn_hp'
+WK2 = '8.2218004e-08*dk2factorn_hp'
+PK2 = '-4.306921e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.31386115
+LVOFF = 8.1825756e-09
+WVOFF = 4.5651731e-07
+PVOFF = -2.3966764e-14
+NFACTOR = 2.25
+ETA0 = 0.29909052
+LETA0 = -7.4992535e-09
+WETA0 = -4.3668614e-07
+PETA0 = 2.1965313e-14
+ETAB = -0.1
+U0 = '(0.03316897*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.6467946e-10*du0factorn_hp'
+WU0 = '-1.5139914e-08*du0factorn_hp'
+PU0 = '7.7524614e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '151310.09*dvsatfactorn_hp'
+LVSAT = '-0.0013233973*dvsatfactorn_hp'
+WVSAT = '-0.077062245*dvsatfactorn_hp'
+PVSAT = '3.8762307e-09*dvsatfactorn_hp'
+A0 = -0.9532925
+LA0 = 1.0293085e-07
+WA0 = 5.7211937e-06
+PA0 = -3.0148447e-13
+AGS = 1.5846684
+LAGS = -2.9408821e-08
+WAGS = -1.7124938e-06
+PAGS = 8.6138438e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.0007665733
+LKETA = 1.4704414e-09
+WKETA = 8.5624707e-08
+PKETA = -4.3069228e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0096580226
+LAIGC = 2.205658e-11
+WAIGC = 1.1481017e-09
+PAIGC = -6.4603723e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.9330834
+LUTE = 2.0439158e-08
+WUTE = 1.1220514e-06
+PUTE = -5.9866295e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.302 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '-0.0046771995+dvth0n302_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0755888e-08+dlvth0n302_hp'
+WVTH0 = '2.2263076e-07+dwvth0n302_hp'
+PVTH0 = '-1.1826551e-14+dpvth0n302_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12638887*dk2factorn_hp'
+LK2 = '-1.217101e-09*dk2factorn_hp'
+WK2 = '3.1829243e-08*dk2factorn_hp'
+PK2 = '-1.8075071e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.004120359
+LCDSCB = -4.2593987e-10
+WCDSCB = -6.6219339e-09
+PCDSCB = 3.9612408e-16
+CDSCD = 0
+CIT = 0
+VOFF = 0.42167672
+LVOFF = -2.9992285e-08
+WVOFF = -2.2753291e-07
+PVOFF = 1.1535857e-14
+NFACTOR = 4.2424415
+LNFACTOR = -9.5836434e-08
+WNFACTOR = -1.8529706e-06
+PNFACTOR = 8.9127883e-14
+ETA0 = -0.18504815
+LETA0 = 1.9560414e-08
+WETA0 = 1.3562822e-08
+PETA0 = -3.2001772e-15
+ETAB = -0.1
+U0 = '(0.025883702*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.2776885e-11*du0factorn_hp'
+WU0 = '-8.3646152e-09*du0factorn_hp'
+PU0 = '4.5211174e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 1.7192396e-27
+LUC = -9.3214894e-35
+WUC = -1.8022838e-33
+PUC = 8.6689852e-41
+EU = 2.9
+VSAT = '22950.012*dvsatfactorn_hp'
+LVSAT = '0.0050992211*dvsatfactorn_hp'
+WVSAT = '0.042312625*dvsatfactorn_hp'
+PVSAT = '-2.0968044e-09*dvsatfactorn_hp'
+A0 = 7.9460662
+LA0 = -3.4927925e-07
+WA0 = -2.5552098e-06
+PA0 = 1.1907093e-13
+AGS = -1.3468919
+LAGS = 1.1804866e-07
+WAGS = 1.0138573e-06
+PAGS = -5.0997022e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.14734462
+LKETA = -5.9024344e-09
+WKETA = -5.0692875e-08
+PKETA = 2.5498516e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.01064482
+LAIGC = -3.1034422e-11
+WAIGC = 2.3037981e-10
+PAIGC = -1.5229091e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.20855508
+LKT1 = 4.2592858e-10
+WKT1 = 8.2352251e-09
+PKT1 = -3.9611358e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.94037047
+LUTE = -3.1144051e-08
+WUTE = 1.9882835e-07
+PUTE = -1.189391e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.402 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.70173723+dvth0n402_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.5875398e-08+dlvth0n402_hp'
+WVTH0 = '-8.2540272e-08+dwvth0n402_hp'
+PVTH0 = '3.9981648e-15+dpvth0n402_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '0.013414104*dk2factorn_hp'
+LK2 = '-8.5500479e-09*dk2factorn_hp'
+WK2 = '-2.8565641e-08*dk2factorn_hp'
+PK2 = '1.3603259e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.012634309
+LCDSCB = 5.8065045e-10
+WCDSCB = 6.1608279e-10
+PCDSCB = -3.8722936e-17
+CDSCD = 0
+CIT = 0
+VOFF = -0.16671947
+LVOFF = -3.1657396e-10
+WVOFF = 2.6654247e-08
+PVOFF = -1.2840507e-15
+NFACTOR = 0.026817282
+LNFACTOR = 1.1156174e-07
+WNFACTOR = -3.1820939e-08
+PNFACTOR = -4.6812655e-16
+ETA0 = -0.25059576
+LETA0 = 1.7997152e-08
+WETA0 = 4.1879388e-08
+PETA0 = -2.5248481e-15
+ETAB = -0.1
+U0 = '(-0.0049056392*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6662935e-09*du0factorn_hp'
+WU0 = '4.9363804e-09*du0factorn_hp'
+PU0 = '-2.3196745e-16*du0factorn_hp'
+UA = -5.0772913e-28
+WUA = 3.1109579e-34
+UB = 1e-19
+UC = -1.5988509e-27
+LUC = 6.0288293e-35
+WUC = -3.6886871e-34
+PUC = 2.0376475e-41
+EU = 2.9
+VSAT = '141294.41*dvsatfactorn_hp'
+LVSAT = '-0.0013636604*dvsatfactorn_hp'
+WVSAT = '-0.008812154*dvsatfactorn_hp'
+PVSAT = '6.9516041e-10*dvsatfactorn_hp'
+A0 = 3.2444518
+LA0 = -1.2526656e-07
+WA0 = -5.2411242e-07
+PA0 = 2.2297447e-14
+AGS = 6.3314525
+LAGS = -3.0535198e-07
+WAGS = -2.3031875e-06
+PAGS = 1.3191206e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.26732763
+LKETA = -1.2723002e-08
+WKETA = -1.0252554e-07
+PKETA = 5.4963367e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.011596986
+LAIGC = -9.7472735e-11
+WAIGC = -1.8095561e-10
+PAIGC = 1.347226e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.18233846
+LKT1 = -8.3508832e-10
+WKT1 = -3.0903535e-09
+PKT1 = 1.4864572e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.39405709
+LUTE = -6.4425837e-08
+WUTE = -3.7179031e-08
+PUTE = 2.4838215e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.502 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.22141426+dvth0n502_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '9.1635818e-09+dlvth0n502_hp'
+WVTH0 = '2.9572171e-09+dwvth0n502_hp'
+PVTH0 = '-4.5877359e-16+dpvth0n502_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12081844*dk2factorn_hp'
+LK2 = '-1.9467782e-09*dk2factorn_hp'
+WK2 = '-4.672248e-09*dk2factorn_hp'
+PK2 = '1.8494393e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.024907457
+LCDSCB = 1.1603279e-09
+WCDSCB = 2.8007031e-09
+PCDSCB = -1.4190552e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.13433234
+LVOFF = -2.1437693e-09
+WVOFF = 2.0889337e-08
+PVOFF = -9.5880991e-16
+NFACTOR = -1.6337108
+LNFACTOR = 1.9545091e-07
+WNFACTOR = 2.6375306e-07
+PNFACTOR = -1.54004e-14
+ETA0 = -0.13586333
+LETA0 = 8.1764453e-09
+WETA0 = 2.1457017e-08
+PETA0 = -7.767623e-16
+ETAB = -0.1
+U0 = '(0.023941758*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.5470566e-11*du0factorn_hp'
+WU0 = '-1.9845636e-10*du0factorn_hp'
+PU0 = '6.1879035e-17*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -7.5296889e-27
+LUC = 3.7479266e-34
+WUC = 6.8682044e-34
+PUC = -3.5605303e-41
+EU = 2.9
+VSAT = '83231.29*dvsatfactorn_hp'
+LVSAT = '0.001634761*dvsatfactorn_hp'
+WVSAT = '0.0015230808*dvsatfactorn_hp'
+PVSAT = '1.614414e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = -7.431269
+LAGS = 4.7650795e-07
+WAGS = 1.4657696e-07
+PAGS = -7.2590115e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.60471347
+LKETA = 3.8935451e-08
+WKETA = 5.2697779e-08
+PKETA = -3.6988678e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0098674576
+LAIGC = 2.1969787e-11
+WAIGC = 1.2690039e-10
+PAIGC = -7.7885087e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21474794
+LKT1 = 7.6323168e-10
+WKT1 = 2.6785339e-09
+PKT1 = -1.3585524e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = 0.16209873
+LUTE = -8.9159824e-08
+WUTE = -1.3617477e-07
+PUTE = 6.8864712e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.602 NMOS
+LMIN = '9.30000000e-08+dlminn_hp'
+LMAX = '9.50000000e-08+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.65975434+dvth0n602_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.5063814e-08+dlvth0n602_hp'
+WVTH0 = '-3.8685091e-08+dwvth0n602_hp'
+PVTH0 = '1.842829e-15+dpvth0n602_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.198*dk2factorn_hp'
+WK2 = '2.66e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.020179787
+LCDSCB = -1.2669748e-09
+WCDSCB = -1.4825851e-09
+PCDSCB = 8.8688235e-17
+CDSCD = 0
+CIT = 0
+VOFF = 0.35360831
+LVOFF = -2.8534437e-08
+WVOFF = -2.5465025e-08
+PVOFF = 1.5483035e-15
+NFACTOR = 6.8167344
+LNFACTOR = -3.0694884e-07
+WNFACTOR = -5.3903924e-07
+PNFACTOR = 3.2327577e-14
+ETA0 = 1.5160089
+LETA0 = -7.185712e-08
+WETA0 = -1.3547085e-07
+PETA0 = 6.8264264e-15
+ETAB = -0.1
+U0 = '(-0.033184423*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6357335e-09*du0factorn_hp'
+WU0 = '5.2285309e-09*du0factorn_hp'
+PU0 = '-9.2045947e-17*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -3e-28
+EU = 2.9
+VSAT = '138704.42*dvsatfactorn_hp'
+LVSAT = '-0.0052945351*dvsatfactorn_hp'
+WVSAT = '-0.0037468666*dvsatfactorn_hp'
+PVSAT = '8.1972453e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = -27.975744
+LAGS = 1.5203697e-06
+WAGS = 2.0983021e-06
+PAGS = -1.0642588e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.49525328
+LKETA = -2.6946417e-08
+WKETA = -5.1799061e-08
+PKETA = 2.5599096e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.014068796
+LAIGC = -2.1008798e-10
+WAIGC = -2.7222678e-10
+PAIGC = 1.4256979e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.14974083
+LKT1 = -2.5339292e-09
+WKT1 = -3.497142e-09
+PKT1 = 1.7737504e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -3.4260384
+LUTE = 1.1629435e-07
+WUTE = 2.0469826e-07
+PUTE = -1.2631675e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = -105938.26
+LAT = 0.0058383929
+WAT = 0.014814135
+PAT = -5.5464732e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.003 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.48470208+dvth0n003_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.2288183e-09+dlvth0n003_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13609769*dk2factorn_hp'
+LK2 = '-2.0612027e-10*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0036867047
+LCDSCB = -3.3917477e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.023561144
+LVOFF = -5.4398798e-09
+NFACTOR = 2.0548833
+LNFACTOR = 1.0306065e-08
+ETA0 = -0.036810608
+LETA0 = 7.98838e-09
+ETAB = -0.07906756
+LETAB = -1.1056515e-09
+U0 = '(0.032081002*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.1562496e-10*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '75322.696*dvsatfactorn_hp'
+LVSAT = '0.0020256704*dvsatfactorn_hp'
+A0 = 4.8116321
+LA0 = -1.9432192e-07
+AGS = 0.84390662
+LAGS = 8.2448523e-09
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.20840581
+LKETA = -1.0587486e-08
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.044417554
+LPDIBLC2 = 2.0985732e-10
+PDIBLCB = 0.21170743
+LPDIBLCB = 1.3980926e-12
+DROUT = 0.56
+PVAG = 0.17434479
+LPVAG = 6.6371079e-09
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.989426
+LPDITSD = -1.9852915e-09
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 7.2195331e-10
+LALPHA0 = 4.1224261e-18
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0099306173
+LAIGC = 8.5262935e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21263439
+LKT1 = 7.6080056e-10
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n003_hp'
+PVTH0 = '0.0+dpvth0n003_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.103 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.48435119+dvth0n103_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.2375751e-09+dlvth0n103_hp'
+WVTH0 = '3.4835409e-09+dwvth0n103_hp'
+PVTH0 = '8.6937303e-17+dpvth0n103_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.16000286*dk2factorn_hp'
+LK2 = '1.3328582e-09*dk2factorn_hp'
+WK2 = '2.3733061e-07*dk2factorn_hp'
+PK2 = '-1.5278978e-14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0064850128
+LCDSCB = -4.8111547e-10
+WCDSCB = -2.7781603e-08
+PCDSCB = 1.4091872e-15
+CDSCD = 0
+CIT = 0
+VOFF = -0.13550586
+LVOFF = 1.1682249e-09
+WVOFF = 1.1113872e-06
+PVOFF = -6.5605264e-14
+NFACTOR = 1.9732292
+LNFACTOR = 1.4619034e-08
+WNFACTOR = 8.1066167e-07
+PNFACTOR = -4.281915e-14
+ETA0 = 0.094242951
+LETA0 = 2.7980962e-10
+WETA0 = -1.3010997e-06
+PETA0 = 7.6530686e-14
+ETAB = -0.070307578
+LETAB = -1.5683538e-09
+WETAB = -8.6969105e-08
+PETAB = 4.5937081e-15
+U0 = '(0.044045306*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.131305e-09*du0factorn_hp'
+WU0 = '-1.1878161e-07*du0factorn_hp'
+PU0 = '7.1052711e-15*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '83251.389*dvsatfactorn_hp'
+LVSAT = '0.0013565017*dvsatfactorn_hp'
+WVSAT = '-0.078716061*dvsatfactorn_hp'
+PVSAT = '6.6435073e-09*dvsatfactorn_hp'
+A0 = 4.3554654
+LA0 = -1.6729423e-07
+WA0 = 4.5288237e-06
+PA0 = -2.6833099e-13
+AGS = 1.5990995
+LAGS = -3.1644437e-08
+WAGS = -7.4975552e-06
+PAGS = 3.9602086e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.28306657
+LKETA = -1.5018226e-08
+WKETA = -7.4123198e-07
+PKETA = 4.3988383e-14
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.042754873
+LPDIBLC2 = 2.9768017e-10
+WPDIBLC2 = 1.6507103e-08
+PPDIBLC2 = -8.7190521e-16
+PDIBLCB = 0.21169635
+LPDIBLCB = 1.983178e-12
+WPDIBLCB = 1.0997214e-10
+PPDIBLCB = -5.8087285e-18
+DROUT = 0.56
+PVAG = 0.12175955
+LPVAG = 9.4146603e-09
+WPVAG = 5.2206627e-07
+PPVAG = -2.757554e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.005155
+LPDITSD = -2.8161128e-09
+WPDITSD = -1.5616044e-07
+PPDITSD = 8.2483945e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 6.8929168e-10
+LALPHA0 = 5.8476135e-18
+WALPHA0 = 3.2426467e-16
+PALPHA0 = -1.712766e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0094293732
+LAIGC = 3.5931263e-11
+WAIGC = 4.976352e-09
+PAIGC = -2.7207654e-16
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21804728
+LKT1 = 1.0791867e-09
+WKT1 = 5.3739169e-08
+PKT1 = -3.1609379e-15
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7888842
+LUTE = 1.9286151e-08
+WUTE = 3.2552347e-06
+PUTE = -1.914729e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.203 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.60223473+dvth0n203_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.2836091e-08+dlvth0n203_hp'
+WVTH0 = '-3.4179734e-07+dwvth0n203_hp'
+PVTH0 = '1.941399e-14+dpvth0n203_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.072839109*dk2factorn_hp'
+LK2 = '-4.2199225e-09*dk2factorn_hp'
+WK2 = '-1.7972026e-08*dk2factorn_hp'
+PK2 = '9.8511641e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = 0.27506951
+LVOFF = -2.2924742e-08
+WVOFF = -9.1188091e-08
+PVOFF = 4.9630356e-15
+NFACTOR = 2.25
+ETA0 = -0.43348194
+LETA0 = 3.1195224e-08
+WETA0 = 2.4460648e-07
+PETA0 = -1.4020563e-14
+ETAB = -0.1
+U0 = '(-0.0027414387*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6321084e-09*du0factorn_hp'
+WU0 = '1.8256766e-08*du0factorn_hp'
+PU0 = '-9.887665e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '50760.919*dvsatfactorn_hp'
+LVSAT = '0.0039876097*dvsatfactorn_hp'
+WVSAT = '0.016448524*dvsatfactorn_hp'
+PVSAT = '-1.0630082e-09*dvsatfactorn_hp'
+A0 = 6.2287891
+LA0 = -2.764267e-07
+WA0 = -9.5814154e-07
+PA0 = 5.1318022e-14
+AGS = -1.2881644
+LAGS = 1.2233421e-07
+WAGS = 9.5924076e-07
+PAGS = -5.4982582e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.00076658087
+LKETA = 1.470441e-09
+WKETA = 8.5624685e-08
+PKETA = -4.3069216e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.01123808
+LAIGC = -6.1402038e-11
+WAIGC = -3.2134969e-10
+PAIGC = 1.3012698e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.65467236
+LUTE = -4.7086515e-08
+WUTE = -6.6871916e-08
+PUTE = 2.9326358e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.303 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '-0.0046773114+dvth0n303_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0755894e-08+dlvth0n303_hp'
+WVTH0 = '2.2263086e-07+dwvth0n303_hp'
+PVTH0 = '-1.1826556e-14+dpvth0n303_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12638906*dk2factorn_hp'
+LK2 = '-1.217091e-09*dk2factorn_hp'
+WK2 = '3.1829429e-08*dk2factorn_hp'
+PK2 = '-1.8075169e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0041203587
+LCDSCB = -4.2593985e-10
+WCDSCB = -6.6219335e-09
+PCDSCB = 3.9612406e-16
+CDSCD = 0
+CIT = 0
+VOFF = 0.42167701
+LVOFF = -2.99923e-08
+WVOFF = -2.2753307e-07
+PVOFF = 1.1535865e-14
+NFACTOR = 4.2424422
+LNFACTOR = -9.5836473e-08
+WNFACTOR = -1.8529713e-06
+PNFACTOR = 8.912792e-14
+ETA0 = -0.18504768
+LETA0 = 1.9560389e-08
+WETA0 = 1.3562622e-08
+PETA0 = -3.2001666e-15
+ETAB = -0.1
+U0 = '(0.025883705*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.2776732e-11*du0factorn_hp'
+WU0 = '-8.3646183e-09*du0factorn_hp'
+PU0 = '4.521119e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 1.7192395e-27
+LUC = -9.3214891e-35
+WUC = -1.8022838e-33
+PUC = 8.6689848e-41
+EU = 2.9
+VSAT = '22950.148*dvsatfactorn_hp'
+LVSAT = '0.0050992138*dvsatfactorn_hp'
+WVSAT = '0.042312541*dvsatfactorn_hp'
+PVSAT = '-2.0968e-09*dvsatfactorn_hp'
+A0 = 7.9460673
+LA0 = -3.4927931e-07
+WA0 = -2.5552102e-06
+PA0 = 1.1907095e-13
+AGS = -1.3468918
+LAGS = 1.1804866e-07
+WAGS = 1.0138572e-06
+PAGS = -5.0997019e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.14734459
+LKETA = -5.9024328e-09
+WKETA = -5.0692862e-08
+PKETA = 2.5498509e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010644826
+LAIGC = -3.103471e-11
+WAIGC = 2.3037651e-10
+PAIGC = -1.5228916e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.20855532
+LKT1 = 4.2594098e-10
+WKT1 = 8.2354433e-09
+PKT1 = -3.9612511e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.94037145
+LUTE = -3.1143999e-08
+WUTE = 1.9882824e-07
+PUTE = -1.1893904e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.403 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.70173736+dvth0n403_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.5875405e-08+dlvth0n403_hp'
+WVTH0 = '-8.2540277e-08+dwvth0n403_hp'
+PVTH0 = '3.998165e-15+dpvth0n403_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '0.013414528*dk2factorn_hp'
+LK2 = '-8.5500703e-09*dk2factorn_hp'
+WK2 = '-2.8565721e-08*dk2factorn_hp'
+PK2 = '1.3603302e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.012634308
+LCDSCB = 5.8065036e-10
+WCDSCB = 6.1608231e-10
+PCDSCB = -3.872291e-17
+CDSCD = 0
+CIT = 0
+VOFF = -0.16671964
+LVOFF = -3.165651e-10
+WVOFF = 2.6654285e-08
+PVOFF = -1.2840527e-15
+NFACTOR = 0.026815164
+LNFACTOR = 1.1156185e-07
+WNFACTOR = -3.182039e-08
+PNFACTOR = -4.6815555e-16
+ETA0 = -0.25059576
+LETA0 = 1.7997152e-08
+WETA0 = 4.1879388e-08
+PETA0 = -2.5248481e-15
+ETAB = -0.1
+U0 = '(-0.004905643*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6662937e-09*du0factorn_hp'
+WU0 = '4.9363802e-09*du0factorn_hp'
+PU0 = '-2.3196744e-16*du0factorn_hp'
+UA = -5.0772913e-28
+WUA = 3.1109579e-34
+UB = 1e-19
+UC = -1.5988508e-27
+LUC = 6.0288285e-35
+WUC = -3.6886875e-34
+PUC = 2.0376477e-41
+EU = 2.9
+VSAT = '141294.41*dvsatfactorn_hp'
+LVSAT = '-0.0013636605*dvsatfactorn_hp'
+WVSAT = '-0.0088121798*dvsatfactorn_hp'
+PVSAT = '6.9516177e-10*dvsatfactorn_hp'
+A0 = 3.244452
+LA0 = -1.2526657e-07
+WA0 = -5.2411246e-07
+PA0 = 2.2297449e-14
+AGS = 6.331454
+LAGS = -3.0535206e-07
+WAGS = -2.3031881e-06
+PAGS = 1.3191209e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.26732764
+LKETA = -1.2723002e-08
+WKETA = -1.0252554e-07
+PKETA = 5.4963369e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.011596975
+LAIGC = -9.7472156e-11
+WAIGC = -1.8095182e-10
+PAIGC = 1.347206e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.182338
+LKT1 = -8.3511262e-10
+WKT1 = -3.0904354e-09
+PKT1 = 1.4865005e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.39405824
+LUTE = -6.4425777e-08
+WUTE = -3.7179069e-08
+PUTE = 2.4838235e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.503 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.22141439+dvth0n503_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '9.1635747e-09+dlvth0n503_hp'
+WVTH0 = '2.9572114e-09+dwvth0n503_hp'
+PVTH0 = '-4.5877329e-16+dpvth0n503_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1208185*dk2factorn_hp'
+LK2 = '-1.9467752e-09*dk2factorn_hp'
+WK2 = '-4.6722427e-09*dk2factorn_hp'
+PK2 = '1.8494365e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.024907457
+LCDSCB = 1.1603279e-09
+WCDSCB = 2.8007029e-09
+PCDSCB = -1.4190551e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.13433224
+LVOFF = -2.1437745e-09
+WVOFF = 2.0889327e-08
+PVOFF = -9.588094e-16
+NFACTOR = -1.6337085
+LNFACTOR = 1.9545079e-07
+WNFACTOR = 2.6375282e-07
+PNFACTOR = -1.5400387e-14
+ETA0 = -0.13586332
+LETA0 = 8.1764449e-09
+WETA0 = 2.1457016e-08
+PETA0 = -7.7676226e-16
+ETAB = -0.1
+U0 = '(0.023941741*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.5471495e-11*du0factorn_hp'
+WU0 = '-1.9845416e-10*du0factorn_hp'
+PU0 = '6.1878919e-17*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -7.529689e-27
+LUC = 3.7479267e-34
+WUC = 6.8682045e-34
+PUC = -3.5605303e-41
+EU = 2.9
+VSAT = '83231.009*dvsatfactorn_hp'
+LVSAT = '0.0016347758*dvsatfactorn_hp'
+WVSAT = '0.0015231055*dvsatfactorn_hp'
+PVSAT = '1.614401e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = -7.4312764
+LAGS = 4.7650834e-07
+WAGS = 1.4657789e-07
+PAGS = -7.2590603e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.60471349
+LKETA = 3.8935452e-08
+WKETA = 5.2697782e-08
+PKETA = -3.698868e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0098674706
+LAIGC = 2.19691e-11
+WAIGC = 1.2689991e-10
+PAIGC = -7.7884835e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21474815
+LKT1 = 7.6324282e-10
+WKT1 = 2.6785714e-09
+PKT1 = -1.3585722e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = 0.16209479
+LUTE = -8.9159616e-08
+WUTE = -1.3617431e-07
+PUTE = 6.886447e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.603 NMOS
+LMIN = '9.50000000e-08+dlminn_hp'
+LMAX = '1.01000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.61792923+dvth0n603_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.2854611e-08+dlvth0n603_hp'
+WVTH0 = '-3.4711698e-08+dwvth0n603_hp'
+PVTH0 = '1.6329544e-15+dpvth0n603_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.18656735*dk2factorn_hp'
+LK2 = '-6.0387243e-10*dk2factorn_hp'
+WK2 = '1.5738985e-09*dk2factorn_hp'
+PK2 = '5.7367881e-17*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.019036528
+LCDSCB = -1.2065879e-09
+WCDSCB = -1.3739757e-09
+PCDSCB = 8.2951488e-17
+CDSCD = 0
+CIT = 0
+VOFF = 0.38037769
+LVOFF = -2.9948395e-08
+WVOFF = -2.8008116e-08
+PVOFF = 1.6826296e-15
+NFACTOR = 6.5134223
+LNFACTOR = -2.9092789e-07
+WNFACTOR = -5.102246e-07
+PNFACTOR = 3.0805588e-14
+ETA0 = 1.4568733
+LETA0 = -6.8733578e-08
+WETA0 = -1.2985296e-07
+PETA0 = 6.5296899e-15
+ETAB = -0.130662
+LETAB = 1.619567e-09
+WETAB = 2.9128903e-09
+PETAB = -1.5385887e-16
+U0 = '(-0.030779682*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.5087152e-09*du0factorn_hp'
+WU0 = '5.000081e-09*du0factorn_hp'
+PU0 = '-7.9979228e-17*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -3e-28
+EU = 2.9
+VSAT = '123920.43*dvsatfactorn_hp'
+LVSAT = '-0.0045136445*dvsatfactorn_hp'
+WVSAT = '-0.0023423892*dvsatfactorn_hp'
+PVSAT = '7.4554003e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = -26.832484
+LAGS = 1.4599828e-06
+WAGS = 1.9896926e-06
+PAGS = -1.0068913e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.43020559
+LKETA = -2.3510598e-08
+WKETA = -4.5619531e-08
+PKETA = 2.2335068e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.054210483
+LPDIBLC2 = -3.0740514e-10
+WPDIBLC2 = -5.5288694e-10
+PPDIBLC2 = 2.9203488e-17
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.4143251
+LPVAG = -6.0386518e-09
+WPVAG = -1.0860885e-08
+PPVAG = 5.7367192e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.896777
+LPDITSD = 2.9084468e-09
+WPDITSD = 5.2310195e-09
+PPDITSD = -2.7630245e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 9.143251e-10
+LALPHA0 = -6.0386518e-18
+WALPHA0 = -1.0860885e-17
+PALPHA0 = 5.7367192e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.014055108
+LAIGC = -2.0936499e-10
+WAIGC = -2.7092567e-10
+PAIGC = 1.4188255e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.14974013
+LKT1 = -2.5339662e-09
+WKT1 = -3.497191e-09
+PKT1 = 1.7737763e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -3.379945
+LUTE = 1.138597e-07
+WUTE = 2.0031948e-07
+PUTE = -1.2400388e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = -87843.155
+LAT = 0.0048826095
+WAT = 0.0130951
+PAT = -4.638479e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.004 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30975798+dvth0n004_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0613935e-09+dlvth0n004_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1165856*dk2factorn_hp'
+LK2 = '-1.3538213e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0066828033
+LCDSCB = 2.7075969e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.060806264
+LVOFF = -3.2491219e-09
+NFACTOR = 1.0792977
+LNFACTOR = 6.769001e-08
+ETA0 = 0.099
+ETAB = 0.025594624
+LETAB = -7.2618812e-09
+U0 = '(0.037443516*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.3104802e-10*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '95951.713*dvsatfactorn_hp'
+LVSAT = '0.00081227167*dvsatfactorn_hp'
+A0 = 1.9682821
+LA0 = -2.7076074e-08
+AGS = 0.063439345
+LAGS = 5.4151937e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.063656065
+LKETA = 5.4151937e-09
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.024552294
+LPDIBLC2 = 1.378332e-09
+PDIBLCB = 0.21157507
+LPDIBLCB = 9.1835784e-12
+DROUT = 0.56
+PVAG = -0.45393117
+LPVAG = 4.35923e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.177367
+LPDITSD = -1.3039978e-08
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.3171967e-10
+LALPHA0 = 2.7075969e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010397764
+LAIGC = -1.8951246e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n004_hp'
+PVTH0 = '0.0+dpvth0n004_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.104 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.23222268+dvth0n104_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '8.5926243e-09+dlvth0n104_hp'
+WVTH0 = '7.6977045e-07+dwvth0n104_hp'
+PVTH0 = '-4.4986059e-14+dpvth0n104_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11520526*dk2factorn_hp'
+LK2 = '-1.3021366e-09*dk2factorn_hp'
+WK2 = '-1.3703944e-08*dk2factorn_hp'
+PK2 = '-5.1312561e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0019174925
+LCDSCB = 1.3119896e-11
+WCDSCB = -4.7310005e-08
+PCDSCB = 2.5578478e-15
+CDSCD = 0
+CIT = 0
+VOFF = 0.02157104
+LVOFF = -8.0710385e-09
+WVOFF = -8.1784187e-07
+PVOFF = 4.7871988e-14
+NFACTOR = 1.5794961
+LNFACTOR = 3.7778415e-08
+WNFACTOR = -4.9659698e-06
+PNFACTOR = 2.9696231e-13
+ETA0 = 0.099
+ETAB = 0.021773373
+LETAB = -6.9845552e-09
+WETAB = 3.7937386e-08
+PETAB = -2.7532917e-15
+U0 = '(0.030879773*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.5690829e-10*du0factorn_hp'
+WU0 = '6.5164843e-08*du0factorn_hp'
+PU0 = '-3.7144593e-15*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 4.119521e-28
+LUC = -3.7094957e-35
+WUC = -6.2611141e-33
+PUC = 3.6827873e-40
+EU = 2.9
+VSAT = '103542.08*dvsatfactorn_hp'
+LVSAT = '0.00016300299*dvsatfactorn_hp'
+WVSAT = '-0.075357206*dvsatfactorn_hp'
+PVSAT = '6.4459395e-09*dvsatfactorn_hp'
+A0 = 2.1327199
+LA0 = -3.6552337e-08
+WA0 = -1.6325385e-06
+PA0 = 9.4080338e-14
+AGS = -0.66523753
+LAGS = 1.0154387e-07
+WAGS = 7.234304e-06
+PAGS = -4.7050709e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.10285004
+LKETA = 7.6813893e-09
+WKETA = 3.8911776e-07
+PKETA = -2.2498789e-14
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.025277604
+LPDIBLC2 = 1.3256931e-09
+WPDIBLC2 = -7.2008854e-09
+PPDIBLC2 = 5.225987e-16
+PDIBLCB = 0.21157995
+LPDIBLCB = 8.8301788e-12
+WPDIBLCB = -4.8431118e-11
+PPDIBLCB = 3.5085512e-18
+DROUT = 0.56
+PVAG = -0.43099253
+LPVAG = 4.1927538e-08
+WPVAG = -2.2773485e-07
+PPVAG = 1.6527761e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.17051
+LPDITSD = -1.2542273e-08
+WPDITSD = 6.8076283e-08
+PPDITSD = -4.9412096e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.4596709e-10
+LALPHA0 = 2.6041966e-17
+WALPHA0 = -1.4144839e-16
+PALPHA0 = 1.0265582e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010728504
+LAIGC = -4.0483589e-11
+WAIGC = -3.2835875e-09
+PAIGC = 2.137731e-16
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.204 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.61614279+dvth0n204_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.3654163e-08+dlvth0n204_hp'
+WVTH0 = '-3.5473156e-07+dwvth0n204_hp'
+PVTH0 = '2.0174781e-14+dpvth0n204_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13278032*dk2factorn_hp'
+LK2 = '-6.9418023e-10*dk2factorn_hp'
+WK2 = '3.7773405e-08*dk2factorn_hp'
+PK2 = '-2.2938299e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.025080711
+LCDSCB = 1.2987874e-09
+WCDSCB = 2.0535061e-08
+PCDSCB = -1.2078723e-15
+CDSCD = 0
+CIT = 0
+VOFF = -0.45987329
+LVOFF = 2.0304594e-08
+WVOFF = 5.9230858e-07
+PVOFF = -3.5240239e-14
+NFACTOR = -1.2166712
+LNFACTOR = 2.039096e-07
+WNFACTOR = 3.2240042e-06
+PNFACTOR = -1.8963593e-13
+ETA0 = 0.22436364
+LETA0 = -7.4992528e-09
+WETA0 = -3.6719009e-07
+PETA0 = 2.1965311e-14
+ETAB = 0.0974045
+LETAB = -1.1611333e-08
+WETAB = -1.8358618e-07
+PETAB = 1.0798539e-14
+U0 = '(0.069987219*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.6457913e-09*du0factorn_hp'
+WU0 = '-4.9380868e-08*du0factorn_hp'
+PU0 = '2.9896791e-15*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.4267711e-27
+LUC = 1.2987874e-34
+WUC = 2.0535061e-33
+PUC = -1.2078723e-40
+EU = 2.9
+VSAT = '82171.75*dvsatfactorn_hp'
+LVSAT = '0.0021400247*dvsatfactorn_hp'
+WVSAT = '-0.012763498*dvsatfactorn_hp'
+PVSAT = '6.5524297e-10*dvsatfactorn_hp'
+A0 = -0.11027305
+LA0 = 9.6436938e-08
+WA0 = 4.9371878e-06
+PA0 = -2.9544525e-13
+AGS = 2.7636694
+LAGS = -1.1599466e-07
+WAGS = -2.8089645e-06
+PAGS = 1.6666325e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.00076658574
+LKETA = 1.4704407e-09
+WKETA = 8.562467e-08
+PKETA = -4.3069208e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.010922432
+LPDIBLC2 = 2.2038788e-09
+WPDIBLC2 = 3.4845415e-08
+PPDIBLC2 = -2.0496073e-15
+PDIBLCB = 0.2114841
+LPDIBLCB = 1.4693419e-11
+WPDIBLCB = 2.323169e-10
+PPDIBLCB = -1.366488e-17
+DROUT = 0.56
+PVAG = -0.88499848
+LPVAG = 6.970161e-08
+WPVAG = 1.1020486e-06
+PPVAG = -6.4822498e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.306297
+LPDITSD = -2.0849188e-08
+WPDITSD = -3.2964545e-07
+PPDITSD = 1.9389745e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 6.3976602e-11
+LALPHA0 = 4.3292896e-17
+WALPHA0 = 6.8450176e-16
+PALPHA0 = -4.0262394e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0090095731
+LAIGC = 6.9678722e-11
+WAIGC = 1.7511598e-09
+PAIGC = -1.0889231e-16
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.8026764
+LUTE = 2.0439084e-08
+WUTE = 1.0007703e-06
+PUTE = -5.9866078e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.304 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '-0.0046764944+dvth0n304_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0755846e-08+dlvth0n304_hp'
+WVTH0 = '2.2263037e-07+dwvth0n304_hp'
+PVTH0 = '-1.1826527e-14+dpvth0n304_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1263886*dk2factorn_hp'
+LK2 = '-1.2171181e-09*dk2factorn_hp'
+WK2 = '3.1829101e-08*dk2factorn_hp'
+PK2 = '-1.8074976e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0041203574
+LCDSCB = -4.2593978e-10
+WCDSCB = -6.6219324e-09
+PCDSCB = 3.96124e-16
+CDSCD = 0
+CIT = 0
+VOFF = 0.42167662
+LVOFF = -2.9992277e-08
+WVOFF = -2.2753284e-07
+PVOFF = 1.1535852e-14
+NFACTOR = 4.2424414
+LNFACTOR = -9.5836421e-08
+WNFACTOR = -1.8529705e-06
+PNFACTOR = 8.9127871e-14
+ETA0 = -0.18504804
+LETA0 = 1.956041e-08
+WETA0 = 1.3562763e-08
+PETA0 = -3.2001749e-15
+ETAB = -0.1
+U0 = '(0.025883768*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.2773025e-11*du0factorn_hp'
+WU0 = '-8.3646586e-09*du0factorn_hp'
+PU0 = '4.5211427e-16*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 1.7192397e-27
+LUC = -9.32149e-35
+WUC = -1.8022839e-33
+PUC = 8.6689857e-41
+EU = 2.9
+VSAT = '22950.005*dvsatfactorn_hp'
+LVSAT = '0.0050992223*dvsatfactorn_hp'
+WVSAT = '0.042312725*dvsatfactorn_hp'
+PVSAT = '-2.0968108e-09*dvsatfactorn_hp'
+A0 = 7.9460706
+LA0 = -3.4927951e-07
+WA0 = -2.5552118e-06
+PA0 = 1.1907105e-13
+AGS = -1.3468914
+LAGS = 1.1804863e-07
+WAGS = 1.0138571e-06
+PAGS = -5.0997009e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.14734457
+LKETA = -5.9024316e-09
+WKETA = -5.0692854e-08
+PKETA = 2.5498505e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.04839062
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.3
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.95184
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 8e-10
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010644818
+LAIGC = -3.1034246e-11
+WAIGC = 2.3038217e-10
+PAIGC = -1.522925e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.20855542
+LKT1 = 4.2594711e-10
+WKT1 = 8.2355403e-09
+PKT1 = -3.9613081e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.94037235
+LUTE = -3.1143946e-08
+WUTE = 1.9882747e-07
+PUTE = -1.189386e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.404 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.6970632+dvth0n404_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.560047e-08+dlvth0n404_hp'
+WVTH0 = '-8.0521173e-08+dwvth0n404_hp'
+PVTH0 = '3.8794013e-15+dpvth0n404_hp'
+K1 = '0.89183943*dk1factorn_hp'
+LK1 = '-1.4107355e-08*dk1factorn_hp'
+WK1 = '-1.0361063e-07*dk1factorn_hp'
+PK1 = '6.0943775e-15*dk1factorn_hp'
+K2 = '-0.10766335*dk2factorn_hp'
+LK2 = '-1.4282693e-09*dk2factorn_hp'
+WK2 = '2.3739795e-08*dk2factorn_hp'
+PK2 = '-1.7162803e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.016960386
+LCDSCB = 8.3511028e-10
+WCDSCB = 2.4849487e-09
+PCDSCB = -1.4864963e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.10917112
+LVOFF = -3.7015689e-09
+WVOFF = 1.7933852e-09
+PVOFF = 1.7826545e-16
+NFACTOR = 0.015752776
+LNFACTOR = 1.1221254e-07
+WNFACTOR = -2.7040997e-08
+PNFACTOR = -7.4927946e-16
+ETA0 = 0.02245313
+LETA0 = 1.9364165e-09
+WETA0 = -7.6077741e-08
+PETA0 = 4.4133902e-15
+ETAB = -0.27255434
+LETAB = 1.0149646e-08
+WETAB = 7.4543476e-08
+PETAB = -4.3846472e-15
+U0 = '(-0.0027979749*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.5423207e-09*du0factorn_hp'
+WU0 = '4.0258545e-09*du0factorn_hp'
+PU0 = '-1.7841032e-16*du0factorn_hp'
+UA = 6.1036353e-27
+LUA = -3.8888046e-34
+WUA = -2.5450137e-33
+PUA = 1.6799636e-40
+UB = 1e-19
+UC = -3.8696163e-27
+LUC = 1.9385471e-34
+WUC = 6.1210187e-34
+PUC = -3.7324215e-41
+EU = 2.9
+VSAT = '175350.31*dvsatfactorn_hp'
+LVSAT = '-0.0033668283*dvsatfactorn_hp'
+WVSAT = '-0.023524205*dvsatfactorn_hp'
+PVSAT = '1.5605231e-09*dvsatfactorn_hp'
+A0 = -4.5726078
+LA0 = 3.3453289e-07
+WA0 = 2.8528573e-06
+PA0 = -1.7633591e-13
+AGS = -0.14660111
+LAGS = 7.5687141e-08
+WAGS = 4.9533168e-07
+PAGS = -3.2696845e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.14199019
+LKETA = 1.1353072e-08
+WKETA = 7.4299761e-08
+PKETA = -4.9045272e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.081142613
+LPDIBLC2 = -1.9264722e-09
+WPDIBLC2 = -1.4148861e-08
+PPDIBLC2 = 8.32236e-16
+PDIBLCB = 0.21195189
+LPDIBLCB = -1.2822156e-11
+WPDIBLCB = -9.4171564e-11
+PPDIBLCB = 5.5391714e-18
+DROUT = 0.56
+PVAG = 0.94337951
+LPVAG = -3.7843583e-08
+WPVAG = -2.7793995e-07
+PPVAG = 1.6348428e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.642001
+LPDITSD = 1.8224722e-08
+WPDITSD = 1.3385039e-07
+PPDITSD = -7.87308e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.4433795e-09
+LALPHA0 = -3.7843583e-17
+WALPHA0 = -2.7793995e-16
+PALPHA0 = 1.6348428e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.012435605
+LAIGC = -1.4680042e-10
+WAIGC = -5.4323804e-10
+PAIGC = 3.4781736e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1823378
+LKT1 = -8.3512464e-10
+WKT1 = -3.0904717e-09
+PKT1 = 1.4865219e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = 0.20726229
+LUTE = -9.979545e-08
+WUTE = -2.9695069e-07
+PUTE = 1.776359e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.504 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.23571724+dvth0n504_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '8.322281e-09+dlvth0n504_hp'
+WVTH0 = '1.5984073e-09+dwvth0n504_hp'
+PVTH0 = '-3.7884844e-16+dpvth0n504_hp'
+K1 = '-0.081966449*dk1factorn_hp'
+LK1 = '4.3171907e-08*dk1factorn_hp'
+WK1 = '6.9726813e-08*dk1factorn_hp'
+PK1 = '-4.1013311e-15*dk1factorn_hp'
+K2 = '0.24970745*dk2factorn_hp'
+LK2 = '-2.3741111e-08*dk2factorn_hp'
+WK2 = '-3.9872208e-08*dk2factorn_hp'
+PK2 = '2.2554056e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011668606
+LCDSCB = 3.8161867e-10
+WCDSCB = 1.5430119e-09
+PCDSCB = -6.7928124e-17
+CDSCD = 0
+CIT = 0
+VOFF = -0.3104438
+LVOFF = 8.2151074e-09
+WVOFF = 3.7619921e-08
+PVOFF = -1.9429029e-15
+NFACTOR = -1.5998523
+LNFACTOR = 1.9345937e-07
+WNFACTOR = 2.605367e-07
+PNFACTOR = -1.5211215e-14
+ETA0 = -0.97145884
+LETA0 = 5.7326173e-08
+WETA0 = 1.0083859e-07
+PETA0 = -5.4459864e-15
+ETAB = 0.42805787
+LETAB = -3.1060364e-08
+WETAB = -5.0165497e-08
+PETAB = 2.9507345e-15
+U0 = '(0.017491637*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.9486661e-10*du0factorn_hp'
+WU0 = '4.1430363e-10*du0factorn_hp'
+PU0 = '2.5836506e-17*du0factorn_hp'
+UA = -1.8992368e-26
+LUA = 1.1900679e-33
+WUA = 1.922075e-33
+PUA = -1.1305645e-40
+UB = 1e-19
+UC = -5.8060028e-28
+LUC = -3.395273e-35
+WUC = 2.6657027e-35
+PUC = 3.2255093e-42
+EU = 2.9
+VSAT = '-20987.033*dvsatfactorn_hp'
+LVSAT = '0.0077648811*dvsatfactorn_hp'
+WVSAT = '0.011423842*dvsatfactorn_hp'
+PVSAT = '-4.209212e-10*dvsatfactorn_hp'
+A0 = 24.222085
+LA0 = -1.4070971e-06
+WA0 = -2.2725981e-06
+PA0 = 1.3367422e-13
+AGS = 12.393134
+LAGS = -6.8956346e-07
+WAGS = -1.7367411e-06
+PAGS = 1.0351776e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.64789768
+LKETA = -3.4743137e-08
+WKETA = -6.630028e-08
+PKETA = 3.300598e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = -0.051838371
+LPDIBLC2 = 5.8954692e-09
+WPDIBLC2 = 9.5217541e-09
+PPDIBLC2 = -5.6006958e-16
+PDIBLCB = 0.2110668
+LPDIBLCB = 3.9238887e-11
+WPDIBLCB = 6.3374605e-11
+PPDIBLCB = -3.7276943e-18
+DROUT = 0.56
+PVAG = -1.6688963
+LPVAG = 1.1581048e-07
+WPVAG = 1.8704515e-07
+PPVAG = -1.1001996e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.900022
+LPDITSD = -5.5772041e-08
+WPDITSD = -9.0077251e-08
+PPDITSD = 5.2983439e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -1.1688963e-09
+LALPHA0 = 1.1581048e-16
+WALPHA0 = 1.8704515e-16
+PALPHA0 = -1.1001996e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0073011145
+LAIGC = 1.7292216e-10
+WAIGC = 3.7070134e-10
+PAIGC = -2.2128884e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21474775
+LKT1 = 7.6321882e-10
+WKT1 = 2.6784988e-09
+PKT1 = -1.3585295e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6781074
+LUTE = 1.9081075e-08
+WUTE = 3.8645111e-08
+PUTE = -3.3964313e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.604 NMOS
+LMIN = '1.01000000e-07+dlminn_hp'
+LMAX = '1.02000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.032369418+dvth0n604_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.1588017e-08+dlvth0n604_hp'
+WVTH0 = '2.0916451e-08+dwvth0n604_hp'
+PVTH0 = '-1.6390934e-15+dpvth0n604_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.026513817*dk2factorn_hp'
+LK2 = '-1.0018221e-08*dk2factorn_hp'
+WK2 = '-1.3631187e-08*dk2factorn_hp'
+PK2 = '9.5173103e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0030310017
+LCDSCB = -2.651428e-10
+WCDSCB = 1.4654916e-10
+PCDSCB = -6.4857841e-18
+CDSCD = 0
+CIT = 0
+VOFF = 0.75514903
+LVOFF = -5.1992445e-08
+WVOFF = -6.3611397e-08
+PVOFF = 3.7768146e-15
+NFACTOR = 2.2670695
+LNFACTOR = -4.115742e-08
+WNFACTOR = -1.0682086e-07
+PNFACTOR = 7.0773799e-15
+ETA0 = 0.62897552
+LETA0 = -2.003663e-08
+WETA0 = -5.1202674e-08
+PETA0 = 1.9034798e-15
+ETAB = -0.55993001
+LETAB = 2.6869111e-08
+WETAB = 4.3693351e-08
+PETAB = -2.5525655e-15
+U0 = '(0.0028865522*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.7153277e-10*du0factorn_hp'
+WU0 = '1.8017867e-09*du0factorn_hp'
+PU0 = '1.0814445e-16*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -3e-28
+EU = 2.9
+VSAT = '-83053.965*dvsatfactorn_hp'
+LVSAT = '0.0076605892*dvsatfactorn_hp'
+WVSAT = '0.0173202*dvsatfactorn_hp'
+PVSAT = '-4.1101348e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = -10.826969
+LAGS = 5.1853833e-07
+WAGS = 4.6916861e-07
+PAGS = -1.1251908e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.4804632
+LKETA = 3.005494e-08
+WKETA = 4.0894004e-08
+PKETA = -2.8552193e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.13568842
+LPDIBLC2 = -5.0999373e-09
+WPDIBLC2 = -8.2932909e-09
+PPDIBLC2 = 4.8449405e-16
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 2.0148768
+LPVAG = -1.001831e-07
+WPVAG = -1.6291329e-07
+PPVAG = 9.5173945e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.125995
+LPDITSD = 4.8245806e-08
+WPDITSD = 7.8455248e-08
+PPDITSD = -4.5833515e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 2.5148768e-09
+LALPHA0 = -1.001831e-16
+WALPHA0 = -1.6291329e-16
+PALPHA0 = 9.5173945e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.013861761
+LAIGC = -1.9799232e-10
+WAIGC = -2.5256011e-10
+PAIGC = 1.3107992e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.14974148
+LKT1 = -2.5338865e-09
+WKT1 = -3.4970962e-09
+PKT1 = 1.7737205e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -2.7346858
+LUTE = 7.5905547e-08
+WUTE = 1.3902006e-07
+PUTE = -8.7947562e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 165487.68
+LAT = -0.01001831
+WAT = -0.010971329
+PAT = 9.5173945e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.005 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.309758+dvth0n005_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0613921e-09+dlvth0n005_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11658607*dk2factorn_hp'
+LK2 = '-1.353793e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0066828027
+LCDSCB = 2.7075965e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.060806357
+LVOFF = -3.2491163e-09
+NFACTOR = 1.0792993
+LNFACTOR = 6.7689913e-08
+ETA0 = 0.099
+ETAB = 0.025594641
+LETAB = -7.2618821e-09
+U0 = '(0.037443574*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.310515e-10*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '95951.644*dvsatfactorn_hp'
+LVSAT = '0.0008122758*dvsatfactorn_hp'
+A0 = 1.9682807
+LA0 = -2.7075991e-08
+AGS = 0.06343947
+LAGS = 5.415193e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.063656053
+LKETA = 5.415193e-09
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.024552251
+LPDIBLC2 = 1.3783345e-09
+PDIBLCB = 0.21157523
+LPDIBLCB = 9.1740311e-12
+DROUT = 0.56
+PVAG = -0.45393125
+LPVAG = 4.3592305e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.177365
+LPDITSD = -1.3039855e-08
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.3171973e-10
+LALPHA0 = 2.7075965e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010397806
+LAIGC = -1.8953758e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n005_hp'
+PVTH0 = '0.0+dpvth0n005_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.105 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.23222275+dvth0n105_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '8.5926198e-09+dlvth0n105_hp'
+WVTH0 = '7.6976994e-07+dwvth0n105_hp'
+PVTH0 = '-4.4986028e-14+dpvth0n105_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11520605*dk2factorn_hp'
+LK2 = '-1.3020898e-09*dk2factorn_hp'
+WK2 = '-1.370087e-08*dk2factorn_hp'
+PK2 = '-5.133095e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0019174903
+LCDSCB = 1.3119766e-11
+WCDSCB = -4.7310021e-08
+PCDSCB = 2.5578488e-15
+CDSCD = 0
+CIT = 0
+VOFF = 0.021570888
+LVOFF = -8.0710294e-09
+WVOFF = -8.1784128e-07
+PVOFF = 4.7871953e-14
+NFACTOR = 1.5794987
+LNFACTOR = 3.7778256e-08
+WNFACTOR = -4.96598e-06
+PNFACTOR = 2.9696292e-13
+ETA0 = 0.099
+ETAB = 0.021773387
+LETAB = -6.9845561e-09
+WETAB = 3.7937413e-08
+PETAB = -2.7532933e-15
+U0 = '(0.030879865*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.5691379e-10*du0factorn_hp'
+WU0 = '6.5164507e-08*du0factorn_hp'
+PU0 = '-3.7144392e-15*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 4.1195223e-28
+LUC = -3.7094964e-35
+WUC = -6.2611154e-33
+PUC = 3.6827881e-40
+EU = 2.9
+VSAT = '103542.06*dvsatfactorn_hp'
+LVSAT = '0.0001630046*dvsatfactorn_hp'
+WVSAT = '-0.075357624*dvsatfactorn_hp'
+PVSAT = '6.4459645e-09*dvsatfactorn_hp'
+A0 = 2.1327181
+LA0 = -3.6552232e-08
+WA0 = -1.6325348e-06
+PA0 = 9.4080114e-14
+AGS = -0.66523736
+LAGS = 1.0154386e-07
+WAGS = 7.2343036e-06
+PAGS = -4.7050707e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.10285002
+LKETA = 7.6813882e-09
+WKETA = 3.8911771e-07
+PKETA = -2.2498786e-14
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.025277538
+LPDIBLC2 = 1.325697e-09
+WPDIBLC2 = -7.2006547e-09
+PPDIBLC2 = 5.225849e-16
+PDIBLCB = 0.21158008
+LPDIBLCB = 8.8225141e-12
+WPDIBLCB = -4.811868e-11
+PPDIBLCB = 3.4898612e-18
+DROUT = 0.56
+PVAG = -0.4309927
+LPVAG = 4.1927548e-08
+WPVAG = -2.2773399e-07
+PPVAG = 1.652771e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.170505
+LPDITSD = -1.2541964e-08
+WPDITSD = 6.8107236e-08
+PPDITSD = -4.9430612e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.4596731e-10
+LALPHA0 = 2.6041953e-17
+WALPHA0 = -1.4144989e-16
+PALPHA0 = 1.0265672e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010728564
+LAIGC = -4.0487198e-11
+WAIGC = -3.2837695e-09
+PAIGC = 2.1378399e-16
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.205 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.49376051+dvth0n205_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.3332548e-09+dlvth0n205_hp'
+WVTH0 = '3.7258503e-09+dwvth0n205_hp'
+PVTH0 = '-1.2681417e-15+dpvth0n205_hp'
+K1 = '0.77006703*dk1factorn_hp'
+LK1 = '-7.0627698e-09*dk1factorn_hp'
+WK1 = '-3.4581833e-07*dk1factorn_hp'
+PK1 = '2.0686853e-14*dk1factorn_hp'
+K2 = '-0.16362472*dk2factorn_hp'
+LK2 = '1.1509317e-09*dk2factorn_hp'
+WK2 = '1.2811743e-07*dk2factorn_hp'
+PK2 = '-7.6982094e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.025080715
+LCDSCB = 1.2987877e-09
+WCDSCB = 2.0535065e-08
+PCDSCB = -1.2078725e-15
+CDSCD = 0
+CIT = 0
+VOFF = -0.26607709
+LVOFF = 8.7117048e-09
+WVOFF = 2.4679646e-08
+PVOFF = -1.2846758e-15
+NFACTOR = 0.47159805
+LNFACTOR = 1.0291733e-07
+WNFACTOR = -1.7209388e-06
+PNFACTOR = 1.0617056e-13
+ETA0 = 0.099
+ETAB = 0.012459087
+LETAB = -6.5298981e-09
+WETAB = 6.5218995e-08
+PETAB = -4.0849864e-15
+U0 = '(0.060495083*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0779717e-09*du0factorn_hp'
+WU0 = '-2.1578466e-08*du0factorn_hp'
+PU0 = '1.3265394e-15*du0factorn_hp'
+UA = -7.3775857e-28
+LUA = 5.6838486e-35
+WUA = 2.7830145e-33
+PUA = -1.6647993e-40
+UB = 1e-19
+UC = -9.952547e-28
+LUC = 4.4245431e-35
+WUC = -2.1394063e-33
+PUC = 1.3003279e-40
+EU = 2.9
+VSAT = '79051.715*dvsatfactorn_hp'
+LVSAT = '0.0023266652*dvsatfactorn_hp'
+WVSAT = '-0.0036254099*dvsatfactorn_hp'
+PVSAT = '1.0860256e-10*dvsatfactorn_hp'
+A0 = 1.5628956
+LA0 = -3.6520106e-09
+WA0 = 3.647538e-08
+PA0 = -2.2846331e-15
+AGS = 1.6386086
+LAGS = -4.8693521e-08
+WAGS = 4.8633863e-07
+PAGS = -3.0461781e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.0063242786
+LKETA = 1.8946162e-09
+WKETA = 1.0639381e-07
+PKETA = -5.5493308e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.027045438
+LPDIBLC2 = 1.2394006e-09
+WPDIBLC2 = -1.2378833e-08
+PPDIBLC2 = 7.753472e-16
+PDIBLCB = 0.21159182
+LPDIBLCB = 8.2493803e-12
+WPDIBLCB = -8.251844e-11
+PPDIBLCB = 5.16857e-18
+DROUT = 0.56
+PVAG = -0.56827877
+LPVAG = 5.0755438e-08
+WPVAG = 1.7437693e-07
+PPVAG = -9.3291794e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.153774
+LPDITSD = -1.1725237e-08
+WPDITSD = 1.1711151e-07
+PPDITSD = -7.335256e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.8069569e-10
+LALPHA0 = 2.4346761e-17
+WALPHA0 = -2.4316932e-16
+PALPHA0 = 1.523089e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0095366459
+LAIGC = 3.8149229e-11
+WAIGC = 2.0735834e-10
+PAIGC = -1.6542107e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.305 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.66261323+dvth0n305_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.9161426e-08+dlvth0n305_hp'
+WVTH0 = '-1.5330718e-07+dwvth0n305_hp'
+PVTH0 = '1.0662057e-14+dpvth0n305_hp'
+K1 = '0.36454829*dk1factorn_hp'
+LK1 = '1.7195361e-08*dk1factorn_hp'
+WK1 = '3.1314095e-08*dk1factorn_hp'
+PK1 = '-1.8732091e-15*dk1factorn_hp'
+K2 = '0.03572953*dk2factorn_hp'
+LK2 = '-1.0915025e-08*dk2factorn_hp'
+WK2 = '-5.7282025e-08*dk2factorn_hp'
+PK2 = '3.5231299e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.29853364
+LVOFF = 1.30907e-08
+WVOFF = 5.4864238e-08
+PVOFF = -5.3571417e-15
+NFACTOR = -3.7563163
+LNFACTOR = 3.8264926e-07
+WNFACTOR = 2.2110215e-06
+PNFACTOR = -1.5398013e-13
+ETA0 = 0.38955333
+LETA0 = -1.4812244e-08
+WETA0 = -2.702146e-07
+PETA0 = 1.3775387e-14
+ETAB = 0.10681426
+LETAB = -1.2371629e-08
+WETAB = -2.2531314e-08
+PETAB = 1.3478232e-15
+U0 = '(0.033102099*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.490275e-10*du0factorn_hp'
+WU0 = '3.8970091e-09*du0factorn_hp'
+PU0 = '-2.8137869e-16*du0factorn_hp'
+UA = 3.0879595e-27
+LUA = -1.7201597e-34
+WUA = -7.7490337e-34
+PUA = 4.635472e-41
+UB = 1e-19
+UC = -5.5137125e-27
+LUC = 3.394603e-34
+WUC = 2.0627595e-33
+PUC = -1.4451704e-40
+EU = 2.9
+VSAT = '21908.413*dvsatfactorn_hp'
+LVSAT = '0.0051615303*dvsatfactorn_hp'
+WVSAT = '0.04951786*dvsatfactorn_hp'
+PVSAT = '-2.527822e-09*dvsatfactorn_hp'
+A0 = -1.2787118
+LA0 = 2.0254697e-07
+WA0 = 2.6791703e-06
+PA0 = -1.9404969e-13
+AGS = 3.169166
+LAGS = -1.5210192e-07
+WAGS = -9.370797e-07
+PAGS = 6.5708029e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.27585359
+LKETA = -1.3589841e-08
+WKETA = -1.5603161e-07
+PKETA = 8.8512146e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.0091368259
+LPDIBLC2 = 2.348162e-09
+WPDIBLC2 = 4.2761765e-09
+PPDIBLC2 = -2.5580088e-16
+PDIBLCB = 0.21147245
+LPDIBLCB = 1.5639986e-11
+WPDIBLCB = 2.8497047e-11
+PPDIBLCB = -1.7046933e-18
+DROUT = 0.56
+PVAG = -0.47110052
+LPVAG = 4.6127233e-08
+WPVAG = 8.4001151e-08
+PPVAG = -5.0249489e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.323199
+LPDITSD = -2.2214677e-08
+WPDITSD = -4.0453416e-08
+PPDITSD = 2.4199234e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 2.8899483e-11
+LALPHA0 = 4.6127233e-17
+WALPHA0 = 8.4001151e-17
+PALPHA0 = -5.0249489e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0098905419
+LAIGC = 1.4086542e-11
+WAIGC = -1.2176497e-10
+PAIGC = 5.8361923e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.19143033
+LKT1 = -5.9847567e-10
+WKT1 = -7.6907917e-09
+PKT1 = 5.5658237e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.405 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.35153453+dvth0n405_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '5.0690545e-09+dlvth0n405_hp'
+WVTH0 = '-1.8921181e-08+dwvth0n405_hp'
+PVTH0 = '1.9448983e-16+dpvth0n405_hp'
+K1 = '0.52500228*dk1factorn_hp'
+LK1 = '7.836843e-09*dk1factorn_hp'
+WK1 = '-3.8002029e-08*dk1factorn_hp'
+PK1 = '2.1696707e-15*dk1factorn_hp'
+K2 = '-0.18209156*dk2factorn_hp'
+LK2 = '3.0240263e-09*dk2factorn_hp'
+WK2 = '3.6816688e-08*dk2factorn_hp'
+PK2 = '-2.4985401e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.22213156
+LVOFF = 3.0557246e-09
+WVOFF = 2.185854e-08
+PVOFF = -1.0220321e-15
+NFACTOR = 2.4049511
+LNFACTOR = -3.0709304e-08
+WNFACTOR = -4.5064598e-07
+PNFACTOR = 2.4590771e-14
+ETA0 = -0.11913503
+LETA0 = 1.040622e-08
+WETA0 = -5.0461227e-08
+PETA0 = 2.8810103e-15
+ETAB = -0.0086304738
+LETAB = -5.6382794e-09
+WETAB = 2.734081e-08
+PETAB = -1.5609838e-15
+U0 = '(0.057720229*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0778783e-09*du0factorn_hp'
+WU0 = '-6.7380233e-09*du0factorn_hp'
+PU0 = '4.6548485e-16*du0factorn_hp'
+UA = 7.90973e-27
+LUA = -4.9692104e-34
+WUA = -2.8579082e-33
+PUA = 1.8671371e-40
+UB = 1e-19
+UC = -9.5365898e-28
+LUC = 1.9422146e-35
+WUC = 9.2816375e-35
+PUC = -6.2605567e-42
+EU = 2.9
+VSAT = '201616.22*dvsatfactorn_hp'
+LVSAT = '-0.0049380553*dvsatfactorn_hp'
+WVSAT = '-0.028115912*dvsatfactorn_hp'
+PVSAT = '1.835199e-09*dvsatfactorn_hp'
+A0 = 0.38579245
+LA0 = 3.7921387e-08
+WA0 = 1.9601044e-06
+PA0 = -1.2293144e-13
+AGS = -0.14001852
+LAGS = 7.529337e-08
+WAGS = 4.92488e-07
+PAGS = -3.2526736e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.33715575
+LKETA = 2.3027876e-08
+WKETA = 1.0878843e-07
+PKETA = -6.9676392e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.03104805
+LPDIBLC2 = 1.0701845e-09
+WPDIBLC2 = -5.1894724e-09
+PPDIBLC2 = 2.9628538e-16
+PDIBLCB = 0.2116184
+LPDIBLCB = 7.1273829e-12
+WPDIBLCB = -3.455237e-11
+PPDIBLCB = 1.9727512e-18
+DROUT = 0.56
+PVAG = -0.040676885
+LPVAG = 2.1022671e-08
+WPVAG = -1.0194186e-07
+PPVAG = 5.820222e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.115912
+LPDITSD = -1.0124633e-08
+WPDITSD = 4.9094381e-08
+PPDITSD = -2.8029755e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.5932311e-10
+LALPHA0 = 2.1022671e-17
+WALPHA0 = -1.0194186e-16
+PALPHA0 = 5.820222e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0097633545
+LAIGC = 1.3053636e-11
+WAIGC = -6.6819993e-11
+PAIGC = 6.282408e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21591376
+LKT1 = 1.1733893e-09
+WKT1 = 2.8860492e-09
+PKT1 = -2.088633e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.505 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.31280569+dvth0n505_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.7108503e-09+dlvth0n505_hp'
+WVTH0 = '-1.2027447e-08+dwvth0n505_hp'
+PVTH0 = '4.3625019e-16+dpvth0n505_hp'
+K1 = '-0.078212319*dk1factorn_hp'
+LK1 = '4.2947334e-08*dk1factorn_hp'
+WK1 = '6.937017e-08*dk1factorn_hp'
+PK1 = '-4.0799968e-15*dk1factorn_hp'
+K2 = '0.37320349*dk2factorn_hp'
+LK2 = '-3.1128645e-08*dk2factorn_hp'
+WK2 = '-6.2025832e-08*dk2factorn_hp'
+PK2 = '3.5806354e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.019822892
+LCDSCB = -1.5022027e-09
+WCDSCB = -4.0624747e-09
+PCDSCB = 2.6739208e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.001481661
+LVOFF = -1.0267008e-08
+WVOFF = -1.7417142e-08
+PVOFF = 1.3494142e-15
+NFACTOR = 0.29355795
+LNFACTOR = 8.0195568e-08
+WNFACTOR = -7.4818005e-08
+PNFACTOR = 4.8497036e-15
+ETA0 = 0.16356913
+LETA0 = -1.05712e-08
+WETA0 = -1.0078257e-07
+PETA0 = 6.6149912e-15
+ETAB = 0.08860389
+LETAB = -1.0754227e-08
+WETAB = 1.0033093e-08
+PETAB = -6.5034515e-16
+U0 = '(-0.0014445479*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.5276292e-09*du0factorn_hp'
+WU0 = '3.793307e-09*du0factorn_hp'
+PU0 = '-1.7629548e-16*du0factorn_hp'
+UA = -1.8888871e-26
+LUA = 1.1838767e-33
+WUA = 1.9122427e-33
+PUA = -1.1246828e-40
+UB = 1e-19
+UC = -5.8355328e-28
+LUC = -3.3776082e-35
+WUC = 2.6937562e-35
+PUC = 3.2087277e-42
+EU = 2.9
+VSAT = '-83773.792*dvsatfactorn_hp'
+LVSAT = '0.011520785*dvsatfactorn_hp'
+WVSAT = '0.02268351*dvsatfactorn_hp'
+PVSAT = '-1.0944746e-09*dvsatfactorn_hp'
+A0 = 24.099705
+LA0 = -1.3997762e-06
+WA0 = -2.2609719e-06
+PA0 = 1.3297874e-13
+AGS = -10.349582
+LAGS = 6.7090578e-07
+WAGS = 2.3097903e-06
+PAGS = -1.3854574e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.64487596
+LKETA = -3.4562377e-08
+WKETA = -6.6013216e-08
+PKETA = 3.2834259e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.012592305
+LPDIBLC2 = 2.0412262e-09
+WPDIBLC2 = -1.9043497e-09
+PPDIBLC2 = 1.2343995e-16
+PDIBLCB = 0.2110699
+LPDIBLCB = 3.9053318e-11
+WPDIBLCB = 6.3079903e-11
+PPDIBLCB = -3.7100652e-18
+DROUT = 0.56
+PVAG = -0.403221
+LPVAG = 4.0097784e-08
+WPVAG = -3.7409005e-08
+PPVAG = 2.4248518e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.290506
+LPDITSD = -1.9310816e-08
+WPDITSD = 1.8016678e-08
+PPDITSD = -1.1678349e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 9.6778996e-11
+LALPHA0 = 4.0097784e-17
+WALPHA0 = -3.7409005e-17
+PALPHA0 = 2.4248518e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0090863206
+LAIGC = 6.6131138e-11
+WAIGC = 5.3692045e-11
+PAIGC = -3.1653875e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.17687711
+LKT1 = -1.5022027e-09
+WKT1 = -4.0624747e-09
+PKT1 = 2.6739208e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -2.4766187
+LUTE = 6.6848021e-08
+WUTE = 1.8078012e-07
+PUTE = -1.1898948e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.605 NMOS
+LMIN = '1.02000000e-07+dlminn_hp'
+LMAX = '1.08000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '-0.21972983+dvth0n605_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.6668594e-08+dlvth0n605_hp'
+WVTH0 = '3.8563427e-08+dwvth0n605_hp'
+PVTH0 = '-2.6947355e-15+dpvth0n605_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.44337221*dk2factorn_hp'
+LK2 = '1.4918248e-08*dk2factorn_hp'
+WK2 = '1.554886e-08*dk2factorn_hp'
+PK2 = '-7.938194e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.10152077
+LCDSCB = 5.9891443e-09
+WCDSCB = 7.4651733e-09
+PCDSCB = -4.4428588e-16
+CDSCD = 0
+CIT = 0
+VOFF = -0.27227833
+LVOFF = 9.4682589e-09
+WVOFF = 8.3085409e-09
+PVOFF = -5.2543612e-16
+NFACTOR = -3.9521621
+LNFACTOR = 3.3087701e-07
+WNFACTOR = 3.285254e-07
+PNFACTOR = -1.8965033e-14
+ETA0 = -3.1227646
+LETA0 = 2.0439246e-07
+WETA0 = 2.1141913e-07
+PETA0 = -1.3806557e-14
+ETAB = 0.55808844
+LETAB = -4.0010752e-08
+WETAB = -3.4567939e-08
+PETAB = 2.1290248e-15
+U0 = '(0.06608934*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.2523235e-09*du0factorn_hp'
+WU0 = '-2.6224123e-09*du0factorn_hp'
+PU0 = '3.7280003e-16*du0factorn_hp'
+UA = 1.24e-27
+UB = 1e-19
+UC = -3e-28
+EU = 2.9
+VSAT = '128744.05*dvsatfactorn_hp'
+LVSAT = '-0.005009168*dvsatfactorn_hp'
+WVSAT = '0.0024943154*dvsatfactorn_hp'
+PVSAT = '4.7587096e-10*dvsatfactorn_hp'
+A0 = 0.3
+AGS = 64.611974
+LAGS = -3.9942192e-06
+WAGS = -4.8115575e-06
+PAGS = 3.0464113e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.48046316
+LKETA = 3.0054938e-08
+WKETA = 4.0894e-08
+PKETA = -2.8552191e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = -0.076519079
+LPDIBLC2 = 7.5943152e-09
+WPDIBLC2 = 6.5612318e-09
+PPDIBLC2 = -4.041035e-16
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = -2.1537226
+LPVAG = 1.4918251e-07
+WPVAG = 1.2888865e-07
+PPVAG = -7.9381974e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 15.133538
+LPDITSD = -7.1845394e-08
+WPDITSD = -6.2071358e-08
+PPDITSD = 3.82295e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -1.6537226e-09
+LALPHA0 = 1.4918251e-16
+WALPHA0 = 1.2888865e-16
+PALPHA0 = -7.9381974e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0079652384
+LAIGC = 1.5473769e-10
+WAIGC = 1.6019485e-10
+PAIGC = -1.158301e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.275472
+LKT1 = 4.987313e-09
+WKT1 = 5.30404e-09
+PKT1 = -3.4911191e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.083624562
+LUTE = -8.2680936e-08
+WUTE = -4.6554317e-08
+PUTE = 2.3063031e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 165487.74
+LAT = -0.010018314
+WAT = -0.010971335
+PAT = 9.5173982e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.006 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30975788+dvth0n006_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0613999e-09+dlvth0n006_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11658591*dk2factorn_hp'
+LK2 = '-1.3538038e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.006682802
+LCDSCB = 2.7075961e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.060806407
+LVOFF = -3.249113e-09
+NFACTOR = 1.0793003
+LNFACTOR = 6.7689844e-08
+ETA0 = 0.099
+ETAB = 0.025594632
+LETAB = -7.2618816e-09
+U0 = '(0.037443554*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.3105014e-10*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '95951.476*dvsatfactorn_hp'
+LVSAT = '0.00081228686*dvsatfactorn_hp'
+A0 = 1.9682802
+LA0 = -2.7075961e-08
+AGS = 0.063439424
+LAGS = 5.4151933e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.063656058
+LKETA = 5.4151933e-09
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.024552246
+LPDIBLC2 = 1.3783348e-09
+PDIBLCB = 0.21157514
+LPDIBLCB = 9.1796159e-12
+DROUT = 0.56
+PVAG = -0.45393111
+LPVAG = 4.3592296e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.177365
+LPDITSD = -1.303988e-08
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.317198e-10
+LALPHA0 = 2.7075961e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010397797
+LAIGC = -1.8953207e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n006_hp'
+PVTH0 = '0.0+dpvth0n006_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.106 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.23222258+dvth0n106_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '8.5926309e-09+dlvth0n106_hp'
+WVTH0 = '7.6977044e-07+dwvth0n106_hp'
+PVTH0 = '-4.4986061e-14+dpvth0n106_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11520583*dk2factorn_hp'
+LK2 = '-1.3021038e-09*dk2factorn_hp'
+WK2 = '-1.3701351e-08*dk2factorn_hp'
+PK2 = '-5.1327785e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0019174897
+LCDSCB = 1.3119722e-11
+WCDSCB = -4.7310021e-08
+PCDSCB = 2.5578488e-15
+CDSCD = 0
+CIT = 0
+VOFF = 0.021570876
+LVOFF = -8.0710286e-09
+WVOFF = -8.1784167e-07
+PVOFF = 4.7871978e-14
+NFACTOR = 1.5795002
+LNFACTOR = 3.7778161e-08
+WNFACTOR = -4.9659841e-06
+PNFACTOR = 2.9696319e-13
+ETA0 = 0.099
+ETAB = 0.021773369
+LETAB = -6.9845549e-09
+WETAB = 3.7937502e-08
+PETAB = -2.7532991e-15
+U0 = '(0.030879834*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.5691177e-10*du0factorn_hp'
+WU0 = '6.5164606e-08*du0factorn_hp'
+PU0 = '-3.7144457e-15*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = 4.1195221e-28
+LUC = -3.7094963e-35
+WUC = -6.2611151e-33
+PUC = 3.6827879e-40
+EU = 2.9
+VSAT = '103541.83*dvsatfactorn_hp'
+LVSAT = '0.00016301955*dvsatfactorn_hp'
+WVSAT = '-0.075357038*dvsatfactorn_hp'
+PVSAT = '6.4459259e-09*dvsatfactorn_hp'
+A0 = 2.1327171
+LA0 = -3.6552167e-08
+WA0 = -1.6325297e-06
+PA0 = 9.4079777e-14
+AGS = -0.66523738
+LAGS = 1.0154386e-07
+WAGS = 7.2343033e-06
+PAGS = -4.7050705e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.10285003
+LKETA = 7.6813886e-09
+WKETA = 3.8911773e-07
+PKETA = -2.2498787e-14
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.025277535
+LPDIBLC2 = 1.3256973e-09
+WPDIBLC2 = -7.2006695e-09
+PPDIBLC2 = 5.2258587e-16
+PDIBLCB = 0.21157998
+LPDIBLCB = 8.8286346e-12
+WPDIBLCB = -4.803787e-11
+PPDIBLCB = 3.4845423e-18
+DROUT = 0.56
+PVAG = -0.43099248
+LPVAG = 4.1927534e-08
+WPVAG = -2.277347e-07
+PPVAG = 1.6527757e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.170502
+LPDITSD = -1.2541775e-08
+WPDITSD = 6.8139518e-08
+PPDITSD = -4.945186e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.4596741e-10
+LALPHA0 = 2.6041946e-17
+WALPHA0 = -1.4145032e-16
+PALPHA0 = 1.02657e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010728548
+LAIGC = -4.048615e-11
+WAIGC = -3.2836946e-09
+PAIGC = 2.1377906e-16
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.206 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.4937605+dvth0n206_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.3332544e-09+dlvth0n206_hp'
+WVTH0 = '3.7258754e-09+dwvth0n206_hp'
+PVTH0 = '-1.2681434e-15+dpvth0n206_hp'
+K1 = '0.77006701*dk1factorn_hp'
+LK1 = '-7.0627683e-09*dk1factorn_hp'
+WK1 = '-3.4581827e-07*dk1factorn_hp'
+PK1 = '2.0686848e-14*dk1factorn_hp'
+K2 = '-0.16362458*dk2factorn_hp'
+LK2 = '1.1509221e-09*dk2factorn_hp'
+WK2 = '1.2811714e-07*dk2factorn_hp'
+PK2 = '-7.6981907e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.025080714
+LCDSCB = 1.2987876e-09
+WCDSCB = 2.0535064e-08
+PCDSCB = -1.2078725e-15
+CDSCD = 0
+CIT = 0
+VOFF = -0.26607731
+LVOFF = 8.7117196e-09
+WVOFF = 2.4679881e-08
+PVOFF = -1.2846913e-15
+NFACTOR = 0.47159781
+LNFACTOR = 1.0291735e-07
+WNFACTOR = -1.720938e-06
+PNFACTOR = 1.0617051e-13
+ETA0 = 0.099
+ETAB = 0.012459109
+LETAB = -6.5298995e-09
+WETAB = 6.5218969e-08
+PETAB = -4.0849847e-15
+U0 = '(0.060495089*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0779721e-09*du0factorn_hp'
+WU0 = '-2.1578475e-08*du0factorn_hp'
+PU0 = '1.32654e-15*du0factorn_hp'
+UA = -7.3775857e-28
+LUA = 5.6838486e-35
+WUA = 2.7830145e-33
+PUA = -1.6647992e-40
+UB = 1e-19
+UC = -9.9525459e-28
+LUC = 4.4245424e-35
+WUC = -2.1394064e-33
+PUC = 1.300328e-40
+EU = 2.9
+VSAT = '79051.686*dvsatfactorn_hp'
+LVSAT = '0.0023266671*dvsatfactorn_hp'
+WVSAT = '-0.0036254056*dvsatfactorn_hp'
+PVSAT = '1.0860228e-10*dvsatfactorn_hp'
+A0 = 1.5628965
+LA0 = -3.6520695e-09
+WA0 = 3.647501e-08
+PA0 = -2.2846088e-15
+AGS = 1.6386085
+LAGS = -4.8693512e-08
+WAGS = 4.8633876e-07
+PAGS = -3.0461789e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.0063242786
+LKETA = 1.8946162e-09
+WKETA = 1.0639381e-07
+PKETA = -5.5493308e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.027045429
+LPDIBLC2 = 1.2394012e-09
+WPDIBLC2 = -1.237883e-08
+PPDIBLC2 = 7.7534703e-16
+PDIBLCB = 0.21159166
+LPDIBLCB = 8.2597985e-12
+WPDIBLCB = -8.2246384e-11
+PPDIBLCB = 5.1506632e-18
+DROUT = 0.56
+PVAG = -0.56827881
+LPVAG = 5.075544e-08
+WPVAG = 1.7437697e-07
+PPVAG = -9.3291818e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.153786
+LPDITSD = -1.1725994e-08
+WPDITSD = 1.1710165e-07
+PPDITSD = -7.3346071e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.8069563e-10
+LALPHA0 = 2.4346764e-17
+WALPHA0 = -2.4316927e-16
+PALPHA0 = 1.5230887e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0095366581
+LAIGC = 3.8148425e-11
+WAIGC = 2.0735084e-10
+PAIGC = -1.6541613e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.306 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.66261337+dvth0n306_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.9161435e-08+dlvth0n306_hp'
+WVTH0 = '-1.5330729e-07+dwvth0n306_hp'
+PVTH0 = '1.0662064e-14+dpvth0n306_hp'
+K1 = '0.36454853*dk1factorn_hp'
+LK1 = '1.7195345e-08*dk1factorn_hp'
+WK1 = '3.1313916e-08*dk1factorn_hp'
+PK1 = '-1.8731974e-15*dk1factorn_hp'
+K2 = '0.035729256*dk2factorn_hp'
+LK2 = '-1.0915007e-08*dk2factorn_hp'
+WK2 = '-5.728192e-08*dk2factorn_hp'
+PK2 = '3.523123e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.003
+CDSCD = 0
+CIT = 0
+VOFF = -0.29853362
+LVOFF = 1.3090699e-08
+WVOFF = 5.4864241e-08
+PVOFF = -5.3571419e-15
+NFACTOR = -3.7563159
+LNFACTOR = 3.8264924e-07
+WNFACTOR = 2.2110217e-06
+PNFACTOR = -1.5398014e-13
+ETA0 = 0.38955333
+LETA0 = -1.4812244e-08
+WETA0 = -2.702146e-07
+PETA0 = 1.3775387e-14
+ETAB = 0.10681425
+LETAB = -1.2371629e-08
+WETAB = -2.2531315e-08
+PETAB = 1.3478233e-15
+U0 = '(0.033102096*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.4902733e-10*du0factorn_hp'
+WU0 = '3.8970081e-09*du0factorn_hp'
+PU0 = '-2.8137862e-16*du0factorn_hp'
+UA = 3.0879594e-27
+LUA = -1.7201596e-34
+WUA = -7.7490329e-34
+PUA = 4.6354714e-41
+UB = 1e-19
+UC = -5.5137126e-27
+LUC = 3.394603e-34
+WUC = 2.0627595e-33
+PUC = -1.4451704e-40
+EU = 2.9
+VSAT = '21908.397*dvsatfactorn_hp'
+LVSAT = '0.0051615314*dvsatfactorn_hp'
+WVSAT = '0.049517853*dvsatfactorn_hp'
+PVSAT = '-2.5278215e-09*dvsatfactorn_hp'
+A0 = -1.2787112
+LA0 = 2.0254694e-07
+WA0 = 2.6791702e-06
+PA0 = -1.9404969e-13
+AGS = 3.169166
+LAGS = -1.5210192e-07
+WAGS = -9.370797e-07
+PAGS = 6.5708029e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.27585359
+LKETA = -1.3589841e-08
+WKETA = -1.560316e-07
+PKETA = 8.8512143e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.0091368032
+LPDIBLC2 = 2.3481635e-09
+WPDIBLC2 = 4.2761915e-09
+PPDIBLC2 = -2.5580187e-16
+PDIBLCB = 0.21147272
+LPDIBLCB = 1.5621971e-11
+WPDIBLCB = 2.8367362e-11
+PPDIBLCB = -1.6961575e-18
+DROUT = 0.56
+PVAG = -0.47110061
+LPVAG = 4.6127239e-08
+WPVAG = 8.4001238e-08
+PPVAG = -5.0249546e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.323201
+LPDITSD = -2.2214859e-08
+WPDITSD = -4.0455138e-08
+PPDITSD = 2.4200367e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 2.889939e-11
+LALPHA0 = 4.6127239e-17
+WALPHA0 = 8.4001238e-17
+PALPHA0 = -5.0249546e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0098905503
+LAIGC = 1.4085991e-11
+WAIGC = -1.2176889e-10
+PAIGC = 5.8364501e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.19143036
+LKT1 = -5.9847381e-10
+WKT1 = -7.6907654e-09
+PKT1 = 5.5658064e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.406 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.27173093+dvth0n406_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.0321728e-08+dlvth0n406_hp'
+WVTH0 = '1.5553925e-08+dwvth0n406_hp'
+PVTH0 = '-2.0746617e-15+dpvth0n406_hp'
+K1 = '0.22069201*dk1factorn_hp'
+LK1 = '2.7866545e-08*dk1factorn_hp'
+WK1 = '9.3459934e-08*dk1factorn_hp'
+PK1 = '-6.4831557e-15*dk1factorn_hp'
+K2 = '-0.021707296*dk2factorn_hp'
+LK2 = '-7.5324663e-09*dk2factorn_hp'
+WK2 = '-3.2469329e-08*dk2factorn_hp'
+PK2 = '2.0618656e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0025696637
+LCDSCB = -3.6659526e-10
+WCDSCB = -2.4060947e-09
+PCDSCB = 1.5836915e-16
+CDSCD = 0.027848318
+LCDSCD = -1.8329763e-09
+WCDSCD = -1.2030474e-08
+PCDSCD = 7.9184577e-16
+CIT = 0
+VOFF = -0.19415419
+LVOFF = 1.2142539e-09
+WVOFF = 9.7723292e-09
+PVOFF = -2.2651771e-16
+NFACTOR = 0.77230566
+LNFACTOR = 7.6751418e-08
+WNFACTOR = 2.5465721e-07
+PNFACTOR = -2.1832285e-14
+ETA0 = -0.38536602
+LETA0 = 2.7929544e-08
+WETA0 = 6.4550561e-08
+PETA0 = -4.6890655e-15
+ETAB = 0.23751361
+LETAB = -2.1839483e-08
+WETAB = -7.8993437e-08
+PETAB = 5.4379364e-15
+U0 = '(0.037025246*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.1573446e-10*du0factorn_hp'
+WU0 = '2.2022076e-09*du0factorn_hp'
+PU0 = '-1.2296114e-16*du0factorn_hp'
+UA = -5.413533e-27
+LUA = 3.8001613e-34
+WUA = 2.8977415e-33
+PUA = -1.9212315e-40
+UB = 1e-19
+UC = 4.5406446e-27
+LUC = -3.4221291e-34
+WUC = -2.2807228e-33
+PUC = 1.4996579e-40
+EU = 2.9
+VSAT = '161756.42*dvsatfactorn_hp'
+LVSAT = '-0.0023144831*dvsatfactorn_hp'
+WVSAT = '-0.010896492*dvsatfactorn_hp'
+PVSAT = '7.0181675e-10*dvsatfactorn_hp'
+A0 = 6.9205535
+LA0 = -3.9219659e-07
+WA0 = -8.6291217e-07
+PA0 = 6.2879517e-14
+AGS = 0.93566231
+LAGS = 4.4920573e-09
+WAGS = 2.7793881e-08
+PAGS = -1.9405688e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.0087137058
+LKETA = 1.4098209e-09
+WKETA = -3.3098532e-08
+PKETA = 2.3713604e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = -0.010507864
+LPDIBLC2 = 3.8053948e-09
+WPDIBLC2 = 1.2762688e-08
+PPDIBLC2 = -8.853258e-16
+PDIBLCB = 0.21134165
+LPDIBLCB = 2.5342572e-11
+WPDIBLCB = 8.4988926e-11
+PPDIBLCB = -5.8954569e-18
+DROUT = 0.56
+PVAG = -0.85700027
+LPVAG = 7.4753076e-08
+WPVAG = 2.5070989e-07
+PPVAG = -1.7391316e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.509041
+LPDITSD = -3.6000363e-08
+WPDITSD = -1.2073774e-07
+PPDITSD = 8.3753747e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 7.5693247e-10
+LALPHA0 = 1.4340231e-18
+WALPHA0 = -2.3050905e-16
+PALPHA0 = 1.4282515e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.009000826
+LAIGC = 6.3243259e-11
+WAIGC = 2.6259201e-10
+PAIGC = -1.539949e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.2159137
+LKT1 = 1.1733857e-09
+WKT1 = 2.8860393e-09
+PKT1 = -2.0886265e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7701161
+LUTE = 2.0346025e-08
+WUTE = 1.3353818e-07
+PUTE = -8.7894827e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.506 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.43042325+dvth0n506_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-4.0307378e-09+dlvth0n506_hp'
+WVTH0 = '-1.2693308e-08+dwvth0n506_hp'
+PVTH0 = '4.8007714e-16+dpvth0n506_hp'
+K1 = '0.85304954*dk1factorn_hp'
+LK1 = '-1.8348321e-08*dk1factorn_hp'
+WK1 = '-1.9099706e-08*dk1factorn_hp'
+PK1 = '1.7430905e-15*dk1factorn_hp'
+K2 = '-0.27263365*dk2factorn_hp'
+LK2 = '1.1380356e-08*dk2factorn_hp'
+WK2 = '1.2195561e-08*dk2factorn_hp'
+PK2 = '-1.3046167e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011862907
+LCDSCB = 5.8335652e-10
+WCDSCB = 1.6290282e-10
+PCDSCB = -1.0722263e-17
+CDSCD = -0.044314537
+LCDSCD = 2.9167829e-09
+WCDSCD = 8.145148e-10
+PCDSCD = -5.3611364e-17
+CIT = 0
+VOFF = -0.16023128
+LVOFF = 1.818921e-10
+WVOFF = 3.7340509e-09
+PVOFF = -4.275732e-17
+NFACTOR = 3.3435221
+LNFACTOR = -1.2055307e-07
+WNFACTOR = -2.0301931e-07
+PNFACTOR = 1.3287913e-14
+ETA0 = -0.048730009
+LETA0 = 3.4023292e-09
+WETA0 = 4.6293508e-09
+PETA0 = -3.2322128e-16
+ETAB = -0.2089214
+LETAB = 8.8288879e-09
+WETAB = 4.7199493e-10
+PETAB = -2.1033643e-17
+U0 = '(0.0082761403*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.8781348e-10*du0factorn_hp'
+WU0 = '7.3195483e-09*du0factorn_hp'
+PU0 = '-4.0839268e-16*du0factorn_hp'
+UA = 2.4113045e-27
+LUA = -2.1810086e-34
+WUA = 1.5049204e-33
+PUA = -8.5658328e-41
+UB = 1e-19
+UC = -1.2132583e-26
+LUC = 7.2638106e-34
+WUC = 6.8711175e-34
+PUC = -4.0243938e-41
+EU = 2.9
+VSAT = '21843.352*dvsatfactorn_hp'
+LVSAT = '0.0045690646*dvsatfactorn_hp'
+WVSAT = '0.014008034*dvsatfactorn_hp'
+PVSAT = '-5.2345474e-10*dvsatfactorn_hp'
+A0 = -0.8685619
+LA0 = 2.4363506e-07
+WA0 = 5.2355038e-07
+PA0 = -5.0298516e-14
+AGS = 4.9612739
+LAGS = -3.3685474e-07
+WAGS = -6.8876497e-07
+PAGS = 5.8819162e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.44205186
+LKETA = 3.6979212e-08
+WKETA = 4.403566e-08
+PKETA = -3.9599912e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.13607982
+LPDIBLC2 = -6.0867223e-09
+WPDIBLC2 = -1.3329921e-08
+PPDIBLC2 = 8.7547105e-16
+PDIBLCB = 0.21191666
+LPDIBLCB = -1.6680471e-11
+WPDIBLCB = -1.7362363e-11
+PPDIBLCB = 1.5846447e-18
+DROUT = 0.56
+PVAG = 0.54470092
+LPVAG = -2.2294437e-08
+WPVAG = 1.2070783e-09
+PPVAG = -1.1685877e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.834015
+LPDITSD = 1.073539e-08
+WPDITSD = -5.8322284e-10
+PPDITSD = 5.6410544e-17
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -7.2788061e-10
+LALPHA0 = 9.437688e-17
+WALPHA0 = 3.3787677e-17
+PALPHA0 = -2.2613138e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010767453
+LAIGC = -4.4521006e-11
+WAIGC = -5.1867615e-11
+PAIGC = 3.7825493e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.5150301
+LUTE = -6.2263739e-08
+WUTE = -8.986714e-08
+PUTE = 5.9150552e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.606 NMOS
+LMIN = '1.08000000e-07+dlminn_hp'
+LMAX = '1.12000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.20058244+dvth0n606_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '9.0036407e-09+dlvth0n606_hp'
+WVTH0 = '9.1415694e-09+dwvth0n606_hp'
+PVTH0 = '-7.5818883e-16+dpvth0n606_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '0.071302395*dk2factorn_hp'
+LK2 = '-1.8957635e-08*dk2factorn_hp'
+WK2 = '-2.0478363e-08*dk2factorn_hp'
+PK2 = '1.5774924e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.052911705
+LCDSCB = 2.7896955e-09
+WCDSCB = 4.0625386e-09
+PCDSCB = -2.2032447e-16
+CDSCD = -0.13581465
+LCDSCD = 8.9393203e-09
+WCDSCD = 9.5070255e-09
+PCDSCD = -6.2575242e-16
+CIT = 0
+VOFF = -0.029478807
+LVOFF = -6.5128054e-09
+WVOFF = -8.6874339e-09
+PVOFF = 5.9323894e-16
+NFACTOR = 2.5096537
+LNFACTOR = -9.4439705e-08
+WNFACTOR = -1.2380181e-07
+PNFACTOR = 1.0807144e-14
+ETA0 = 0.28697544
+LETA0 = -2.0036625e-08
+WETA0 = -2.7262667e-08
+PETA0 = 1.9034794e-15
+ETAB = -0.95495158
+LETAB = 5.9577542e-08
+WETAB = 7.1344862e-08
+PETAB = -4.8421558e-15
+U0 = '(0.24407756*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.5967508e-08*du0factorn_hp'
+WU0 = '-1.5081586e-08*du0factorn_hp'
+PU0 = '1.1928629e-15*du0factorn_hp'
+UA = 6.5887772e-26
+LUA = -4.2551164e-33
+WUA = -4.525344e-33
+PUA = 2.9785815e-40
+UB = 1e-19
+UC = -1.7779346e-26
+LUC = 1.1504905e-33
+WUC = 1.2235542e-33
+PUC = -8.0534338e-41
+EU = 2.9
+VSAT = '183069.77*dvsatfactorn_hp'
+LVSAT = '-0.0085848871*dvsatfactorn_hp'
+WVSAT = '-0.0013084758*dvsatfactorn_hp'
+PVSAT = '7.2617067e-10*dvsatfactorn_hp'
+A0 = 16.80148
+LA0 = -1.0861274e-06
+WA0 = -1.1551036e-06
+PA0 = 7.6028918e-14
+AGS = 2.8510122
+LAGS = 7.0887292e-08
+WAGS = -4.8829012e-07
+PAGS = 2.0083669e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.20883384
+LKETA = 1.2176296e-08
+WKETA = 2.1879948e-08
+PKETA = -1.6037141e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = -0.064289347
+LPDIBLC2 = 6.7893542e-09
+WPDIBLC2 = 5.7051505e-09
+PPDIBLC2 = -3.4775623e-16
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 2.9930237
+LPVAG = -1.8957633e-07
+WPVAG = -2.3138358e-07
+PPVAG = 1.5774921e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 12.654912
+LPDITSD = 9.1297772e-08
+WPDITSD = 1.1143161e-07
+PPDITSD = -7.5970157e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -1.9395622e-09
+LALPHA0 = 1.6799647e-16
+WALPHA0 = 1.4889743e-16
+PALPHA0 = -9.2551753e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010131148
+LAIGC = 1.2177525e-11
+WAIGC = 8.5813834e-12
+PAIGC = -1.603811e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -3.455479
+LUTE = 1.3925452e-07
+WUTE = 1.894755e-07
+PUTE = -1.3229179e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 165487.71
+LAT = -0.010018312
+WAT = -0.010971332
+PAT = 9.517396e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.007 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30975804+dvth0n007_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.061389e-09+dlvth0n007_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11658601*dk2factorn_hp'
+LK2 = '-1.3537963e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0066828031
+LCDSCB = 2.7075968e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.060806393
+LVOFF = -3.249114e-09
+NFACTOR = 1.0792988
+LNFACTOR = 6.7689955e-08
+ETA0 = 0.099
+ETAB = 0.025594641
+LETAB = -7.2618822e-09
+U0 = '(0.037443576*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.3105169e-10*du0factorn_hp'
+UA = 2.124e-28
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '95951.645*dvsatfactorn_hp'
+LVSAT = '0.00081227503*dvsatfactorn_hp'
+A0 = 1.9682797
+LA0 = -2.7075927e-08
+AGS = 0.063439571
+LAGS = 5.4151923e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.063656043
+LKETA = 5.4151923e-09
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.024552254
+LPDIBLC2 = 1.3783343e-09
+PDIBLCB = 0.21157508
+LPDIBLCB = 9.1842058e-12
+DROUT = 0.56
+PVAG = -0.45393125
+LPVAG = 4.3592306e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.177362
+LPDITSD = -1.303963e-08
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.3171969e-10
+LALPHA0 = 2.7075968e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010397787
+LAIGC = -1.8952483e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n007_hp'
+PVTH0 = '0.0+dpvth0n007_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.107 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.2338551+dvth0n107_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '8.4786485e-09+dlvth0n107_hp'
+WVTH0 = '7.5356436e-07+dwvth0n107_hp'
+PVTH0 = '-4.3854552e-14+dpvth0n107_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11492365*dk2factorn_hp'
+LK2 = '-1.321806e-09*dk2factorn_hp'
+WK2 = '-1.6503957e-08*dk2factorn_hp'
+PK2 = '-3.1759991e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0014648894
+LCDSCB = -1.8480832e-11
+WCDSCB = -5.1803447e-08
+PCDSCB = 2.8715798e-15
+CDSCD = 0.00040129513
+LCDSCD = -2.8018426e-11
+WCDSCD = -3.984058e-09
+PCDSCD = 2.7816693e-16
+CIT = 0
+VOFF = 0.020080108
+LVOFF = -7.9669432e-09
+WVOFF = -8.0304118e-07
+PVOFF = 4.6838608e-14
+NFACTOR = 1.5697257
+LNFACTOR = 3.8460614e-08
+WNFACTOR = -4.868959e-06
+PNFACTOR = 2.901889e-13
+ETA0 = 0.10297282
+LETA0 = -2.7738221e-10
+WETA0 = -3.9442145e-08
+PETA0 = 2.7538506e-15
+ETAB = 0.022749759
+LETAB = -7.0527264e-09
+WETAB = 2.824399e-08
+PETAB = -2.0764982e-15
+U0 = '(0.031019892*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.6669064e-10*du0factorn_hp'
+WU0 = '6.3774327e-08*du0factorn_hp'
+PU0 = '-3.6173765e-15*du0factorn_hp'
+UA = 1.6024766e-28
+LUA = 3.6412765e-36
+WUA = 5.1776845e-34
+PUA = -3.6150593e-41
+UB = 1e-19
+UC = 4.1306985e-28
+LUC = -3.7172997e-35
+WUC = -6.2722111e-33
+PUC = 3.6905351e-40
+EU = 2.9
+VSAT = '103692.22*dvsatfactorn_hp'
+LVSAT = '0.00015251965*dvsatfactorn_hp'
+WVSAT = '-0.076848379*dvsatfactorn_hp'
+PVSAT = '6.5500513e-09*dvsatfactorn_hp'
+A0 = 2.1332631
+LA0 = -3.6590289e-08
+WA0 = -1.6379553e-06
+PA0 = 9.4458593e-14
+AGS = -0.65795642
+LAGS = 1.010355e-07
+WAGS = 7.1620194e-06
+PAGS = -4.6546018e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.10285001
+LKETA = 7.6813872e-09
+WKETA = 3.8911767e-07
+PKETA = -2.2498783e-14
+DWG = 0
+DWB = 0
+PCLM = 0.67608674
+LPCLM = 2.2194141e-09
+WPCLM = 3.1558785e-07
+PPCLM = -2.2034344e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.0258266
+LPDIBLC2 = 1.2873616e-09
+WPDIBLC2 = -1.2651701e-08
+PPDIBLC2 = 9.0317689e-16
+PDIBLCB = 0.21606109
+LPDIBLCB = -3.0404226e-10
+WPDIBLCB = -4.4537121e-08
+PPDIBLCB = 3.1097123e-15
+DROUT = 0.56
+PVAG = -0.45134043
+LPVAG = 4.3348227e-08
+WPVAG = -2.5721746e-08
+PPVAG = 2.4232123e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.172252
+LPDITSD = -1.266399e-08
+WPDITSD = 5.0725641e-08
+PPDITSD = -3.7293492e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.5436566e-10
+LALPHA0 = 2.545558e-17
+WALPHA0 = -2.2482919e-16
+PALPHA0 = 1.6087213e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010722124
+LAIGC = -4.0037646e-11
+WAIGC = -3.2200229e-09
+PAIGC = 2.093335e-16
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.207 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.51762939+dvth0n207_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-7.9997802e-09+dlvth0n207_hp'
+WVTH0 = '-7.7610542e-08+dwvth0n207_hp'
+PVTH0 = '4.4107652e-15+dpvth0n207_hp'
+K1 = '0.61234443*dk1factorn_hp'
+LK1 = '3.9494218e-09*dk1factorn_hp'
+WK1 = '1.1615115e-07*dk1factorn_hp'
+PK1 = '-1.1567856e-14*dk1factorn_hp'
+K2 = '-0.08183074*dk2factorn_hp'
+LK2 = '-4.5599236e-09*dk2factorn_hp'
+WK2 = '-1.1343309e-07*dk2factorn_hp'
+PK2 = '9.1668464e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.012851758
+LCDSCB = 4.4496191e-10
+WCDSCB = -1.8451308e-08
+PCDSCB = 1.514156e-15
+CDSCD = 0.016075835
+LCDSCD = -1.1224148e-09
+WCDSCD = -4.9894786e-08
+PCDSCD = 3.483654e-15
+CIT = 0
+VOFF = -0.2618475
+LVOFF = 8.4163938e-09
+WVOFF = 2.2724776e-08
+PVOFF = -1.1481858e-15
+NFACTOR = -0.78805481
+LNFACTOR = 1.908663e-07
+WNFACTOR = 2.0369802e-06
+PNFACTOR = -1.5620734e-13
+ETA0 = 0.25815078
+LETA0 = -1.1111907e-08
+WETA0 = -4.9395839e-07
+PETA0 = 3.4488175e-14
+ETAB = 0.13959466
+LETAB = -1.5406504e-08
+WETAB = -3.1399474e-07
+PETAB = 2.2391716e-14
+U0 = '(0.050866787*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.4057241e-09*du0factorn_hp'
+WU0 = '5.6427733e-09*du0factorn_hp'
+PU0 = '-5.7404754e-16*du0factorn_hp'
+UA = -2.4317261e-27
+LUA = 1.751113e-34
+WUA = 8.1096596e-33
+PUA = -5.3838629e-40
+UB = 1e-19
+UC = 2.2773538e-27
+LUC = -1.8424809e-34
+WUC = -1.1732699e-32
+PUC = 7.9983647e-40
+EU = 2.9
+VSAT = '88101.968*dvsatfactorn_hp'
+LVSAT = '0.0016947764*dvsatfactorn_hp'
+WVSAT = '-0.031184545*dvsatfactorn_hp'
+PVSAT = '2.0327814e-09*dvsatfactorn_hp'
+A0 = 1.598226
+LA0 = -6.1187756e-09
+WA0 = -7.0831459e-08
+PA0 = 5.2075289e-15
+AGS = 2.1096937
+LAGS = -8.1584677e-08
+WAGS = -9.4442769e-07
+PAGS = 6.9434324e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.088428048
+LKETA = -4.7209912e-09
+WKETA = -1.7113575e-07
+PKETA = 1.3827783e-14
+DWG = 0
+DWB = 0
+PCLM = -0.56553353
+LPCLM = 8.8909342e-08
+WPCLM = 3.9522936e-06
+PPCLM = -2.7594914e-13
+PDIBLC1 = 0
+PDIBLC2 = 0.053214061
+LPDIBLC2 = -5.8769266e-10
+WPDIBLC2 = -9.2869574e-08
+PPDIBLC2 = 6.3952107e-15
+PDIBLCB = 0.56588782
+LPDIBLCB = -2.4728698e-08
+WPDIBLCB = -1.0691796e-06
+PPDIBLCB = 7.4649528e-14
+DROUT = 0.56
+PVAG = -0.92013348
+LPVAG = 7.5321933e-08
+WPVAG = 1.3473731e-06
+PPVAG = -9.1227773e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.351401
+LPDITSD = -2.5523478e-08
+WPDITSD = -4.739997e-07
+PPDITSD = 3.3936089e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 6.2742842e-10
+LALPHA0 = 7.1198811e-18
+WALPHA0 = -1.02463e-15
+PALPHA0 = 6.9792476e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0093125911
+LAIGC = 5.3792787e-11
+WAIGC = 9.0849988e-10
+PAIGC = -6.5495839e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.307 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.52200197+dvth0n307_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-9.3439469e-09+dlvth0n307_hp'
+WVTH0 = '-8.1677038e-08+dwvth0n307_hp'
+PVTH0 = '5.6608403e-15+dpvth0n307_hp'
+K1 = '0.90578636*dk1factorn_hp'
+LK1 = '-2.059388e-08*dk1factorn_hp'
+WK1 = '-1.5674984e-07*dk1factorn_hp'
+PK1 = '1.1257414e-14*dk1factorn_hp'
+K2 = '-0.24736642*dk2factorn_hp'
+LK2 = '8.8507339e-09*dk2factorn_hp'
+WK2 = '4.0515102e-08*dk2factorn_hp'
+PK2 = '-3.305065e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.049129816
+LCDSCB = 3.2207837e-09
+WCDSCB = 1.5287285e-08
+PCDSCB = -1.0673583e-15
+CDSCD = -0.058376349
+LCDSCD = 4.0758367e-09
+WCDSCD = 1.9345745e-08
+PCDSCD = -1.3507199e-15
+CIT = 0
+VOFF = -0.29888429
+LVOFF = 1.3115183e-08
+WVOFF = 5.7168992e-08
+PVOFF = -5.5180596e-15
+NFACTOR = 1.6038491
+LNFACTOR = 8.402517e-09
+WNFACTOR = -1.874904e-07
+PNFACTOR = 1.3483974e-14
+ETA0 = -0.36873653
+LETA0 = 3.8131555e-08
+WETA0 = 8.904681e-08
+PETA0 = -1.1308245e-14
+ETAB = -0.33962025
+LETAB = 1.8798428e-08
+WETAB = 1.3167513e-07
+PETAB = -9.4188706e-15
+U0 = '(0.067023552*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.7174234e-09*du0factorn_hp'
+WU0 = '-9.3830184e-09*du0factorn_hp'
+PU0 = '6.4583283e-16*du0factorn_hp'
+UA = 8.9606877e-27
+LUA = -5.8204985e-34
+WUA = -2.4852852e-33
+PUA = 1.6577358e-40
+UB = 1e-19
+UC = -1.4065769e-26
+LUC = 9.3656486e-34
+WUC = 3.4664051e-33
+PUC = -2.4251957e-40
+EU = 2.9
+VSAT = '11984.432*dvsatfactorn_hp'
+LVSAT = '0.0058544226*dvsatfactorn_hp'
+WVSAT = '0.039604764*dvsatfactorn_hp'
+PVSAT = '-1.8356896e-09*dvsatfactorn_hp'
+A0 = -0.50932918
+LA0 = 1.4882868e-07
+WA0 = 1.8891949e-06
+PA0 = -1.3889361e-13
+AGS = 1.1758783
+LAGS = -1.2930575e-08
+WAGS = -7.5979439e-08
+PAGS = 5.5860083e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.083019162
+LKETA = 1.1466654e-08
+WKETA = -1.1689846e-08
+PKETA = -1.226727e-15
+DWG = 0
+DWB = 0
+PCLM = 6.266156
+LPCLM = -3.8807922e-07
+WPCLM = -2.4011777e-06
+PPCLM = 1.6765022e-13
+PDIBLC1 = 0
+PDIBLC2 = -0.11616755
+LPDIBLC2 = 1.1096913e-08
+WPDIBLC2 = 6.4655321e-08
+PPDIBLC2 = -4.4714727e-15
+PDIBLCB = -1.2737553
+LPDIBLCB = 1.0371424e-07
+WPDIBLCB = 6.4168852e-07
+PPDIBLCB = -4.4802408e-14
+DROUT = 0.56
+PVAG = 0.98079227
+LPVAG = -5.5243922e-08
+WPVAG = -4.2048783e-07
+PPVAG = 3.0198472e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.623978
+LPDITSD = 2.6604929e-08
+WPDITSD = 2.0250341e-07
+PPDITSD = -1.4543329e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.5426216e-10
+LALPHA0 = 1.0778958e-16
+WALPHA0 = 3.5334223e-16
+PALPHA0 = -2.3830343e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010623926
+LAIGC = -3.7118322e-11
+WAIGC = -3.1104191e-10
+PAIGC = 1.9051493e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.19400067
+LKT1 = -4.1901481e-10
+WKT1 = -5.3003777e-09
+PKT1 = 3.8968377e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5919002
+LUTE = 9.1394498e-09
+WUTE = 1.2173716e-07
+PUTE = -8.4996883e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.407 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30999654+dvth0n407_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '7.6500226e-09+dlvth0n407_hp'
+WVTH0 = '9.9093075e-09+dwvth0n407_hp'
+PVTH0 = '-1.6805545e-15+dpvth0n407_hp'
+K1 = '0.38364502*dk1factorn_hp'
+LK1 = '1.6489166e-08*dk1factorn_hp'
+WK1 = '6.8815216e-08*dk1factorn_hp'
+PK1 = '-4.7624614e-15*dk1factorn_hp'
+K2 = '-0.10907086*dk2factorn_hp'
+LK2 = '-1.4327421e-09*dk2factorn_hp'
+WK2 = '-1.9228582e-08*dk2factorn_hp'
+PK2 = '1.1373966e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.015423431
+LCDSCB = 8.8968259e-10
+WCDSCB = 7.2612691e-10
+PCDSCB = -6.032256e-17
+CDSCD = 0.0061156713
+LCDSCD = -3.156029e-10
+WCDSCD = -8.5148076e-09
+PCDSCD = 5.4638197e-16
+CIT = 0
+VOFF = -0.18401423
+LVOFF = 5.0628161e-10
+WVOFF = 7.5451249e-09
+PVOFF = -7.1014313e-17
+NFACTOR = 0.35373129
+LNFACTOR = 1.0597628e-07
+WNFACTOR = 3.5256048e-07
+PNFACTOR = -2.8667892e-14
+ETA0 = -0.27656446
+LETA0 = 2.0333019e-08
+WETA0 = 4.9228474e-08
+PETA0 = -3.6192774e-15
+ETAB = 0.099044487
+LETAB = -1.2171569e-08
+WETAB = -5.7828037e-08
+PETAB = 3.9601681e-15
+U0 = '(0.041349361*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.0176442e-09*du0factorn_hp'
+WU0 = '1.7082323e-09*du0factorn_hp'
+PU0 = '-8.8471788e-17*du0factorn_hp'
+UA = -2.8784226e-27
+LUA = 2.0301472e-34
+WUA = 2.6292104e-33
+PUA = -1.7337431e-40
+UB = 1e-19
+UC = -4.2028606e-27
+LUC = 2.6825861e-34
+WUC = -7.9437122e-34
+PUC = 4.6188725e-41
+EU = 2.9
+VSAT = '103327.35*dvsatfactorn_hp'
+LVSAT = '0.0017650344*dvsatfactorn_hp'
+WVSAT = '0.00014462341*dvsatfactorn_hp'
+PVSAT = '-6.9073894e-11*dvsatfactorn_hp'
+A0 = 5.5098215
+LA0 = -2.9369927e-07
+WA0 = -7.1107822e-07
+PA0 = 5.2278471e-14
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.03282211
+LKETA = 3.0930697e-09
+WKETA = -3.3374973e-08
+PKETA = 2.3906615e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.011744628
+LPDIBLC2 = 2.2517258e-09
+WPDIBLC2 = 9.3972616e-09
+PPDIBLC2 = -6.5035175e-16
+PDIBLCB = 0.21148992
+LPDIBLCB = 1.4990397e-11
+WPDIBLCB = 6.2571089e-11
+PPDIBLCB = -4.3302435e-18
+DROUT = 0.56
+PVAG = -0.41987306
+LPVAG = 4.4232854e-08
+WPVAG = 1.8459959e-07
+PPVAG = -1.2775495e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.298529
+LPDITSD = -2.1302411e-08
+WPDITSD = -8.890255e-08
+PPDITSD = 6.1526418e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.2475397e-10
+LALPHA0 = 3.1608726e-17
+WALPHA0 = -1.5599274e-16
+PALPHA0 = 9.0797856e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0094601211
+LAIGC = 3.1175278e-11
+WAIGC = 1.9172196e-10
+PAIGC = -1.0451343e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.21087428
+LKT1 = 8.2153297e-10
+WKT1 = 1.9890216e-09
+PKT1 = -1.4623287e-16
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5288851
+LUTE = 3.5032752e-09
+WUTE = 9.4514661e-08
+PUTE = -6.0648609e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.507 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.44702006+dvth0n507_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.1895269e-09+dlvth0n507_hp'
+WVTH0 = '-1.4480879e-08+dwvth0n507_hp'
+PVTH0 = '6.0488533e-16+dpvth0n507_hp'
+K1 = '0.90559072*dk1factorn_hp'
+LK1 = '-2.2016746e-08*dk1factorn_hp'
+WK1 = '-2.4091119e-08*dk1factorn_hp'
+PK1 = '2.0915909e-15*dk1factorn_hp'
+K2 = '-0.30630856*dk2factorn_hp'
+LK2 = '1.3731538e-08*dk2factorn_hp'
+WK2 = '1.5879729e-08*dk2factorn_hp'
+PK2 = '-1.5618453e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011544098
+LCDSCB = 5.6109726e-10
+WCDSCB = 3.5605587e-11
+PCDSCB = -1.8343708e-18
+CDSCD = -0.042720477
+LCDSCD = 2.8054856e-09
+WCDSCD = 1.7802676e-10
+PCDSCD = -9.1717694e-18
+CIT = 0
+VOFF = -0.16598507
+LVOFF = 5.8362196e-10
+WVOFF = 4.3359354e-09
+PVOFF = -8.4780896e-17
+NFACTOR = 3.6734112
+LNFACTOR = -1.4358593e-07
+WNFACTOR = -2.3834254e-07
+PNFACTOR = 1.5754181e-14
+ETA0 = 0
+ETAB = -0.2294916
+LETAB = 1.0265099e-08
+WETAB = 6.5138651e-10
+PETAB = -3.3558763e-17
+U0 = '(0.0031242316*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.2475197e-09*du0factorn_hp'
+WU0 = '8.5123053e-09*du0factorn_hp'
+PU0 = '-4.9167097e-16*du0factorn_hp'
+UA = 1.8309857e-27
+LUA = -1.77583e-34
+WUA = 1.7909357e-33
+PUA = -1.0562792e-40
+UB = 1e-19
+UC = -1.2223741e-26
+LUC = 7.3274574e-34
+WUC = 6.3334557e-34
+PUC = -3.6489983e-41
+EU = 2.9
+VSAT = '27225.694*dvsatfactorn_hp'
+LVSAT = '0.0041932694*dvsatfactorn_hp'
+WVSAT = '0.013690718*dvsatfactorn_hp'
+PVSAT = '-5.0129973e-10*dvsatfactorn_hp'
+A0 = -2.7747093
+LA0 = 3.7672227e-07
+WA0 = 7.6356826e-07
+PA0 = -6.7056564e-14
+AGS = 5.4656656
+LAGS = -3.7207137e-07
+WAGS = -7.9488847e-07
+PAGS = 6.6228705e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.50877283
+LKETA = 4.163767e-08
+WKETA = 5.1344256e-08
+PKETA = -4.4702773e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.15102724
+LPDIBLC2 = -7.1303512e-09
+WPDIBLC2 = -1.5395044e-08
+PPDIBLC2 = 1.019658e-15
+PDIBLCB = 0.21196454
+LPDIBLCB = -2.0023528e-11
+WPDIBLCB = -2.1911065e-11
+PPDIBLCB = 1.9022351e-18
+DROUT = 0.56
+PVAG = 0.62720499
+LPVAG = -2.8054871e-08
+WPVAG = -1.7802996e-09
+PPVAG = 9.1719955e-17
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.794266
+LPDITSD = 1.3510708e-08
+WPDITSD = 8.562495e-10
+PPDITSD = -4.4093415e-17
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -5.816141e-10
+LALPHA0 = 8.4164551e-17
+WALPHA0 = 5.3407794e-18
+PALPHA0 = -2.7515139e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010886905
+LAIGC = -5.2861134e-11
+WAIGC = -6.2245573e-11
+PAIGC = 4.5071384e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.46785413
+LUTE = -6.5557565e-08
+WUTE = -9.4348858e-08
+PUTE = 6.2279687e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.607 NMOS
+LMIN = '1.12000000e-07+dlminn_hp'
+LMAX = '1.15700000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.50762787+dvth0n607_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.2434272e-08+dlvth0n607_hp'
+WVTH0 = '-2.0238621e-08+dwvth0n607_hp'
+PVTH0 = '1.2931361e-15+dpvth0n607_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '0.0077633186*dk2factorn_hp'
+LK2 = '-1.4521337e-08*dk2factorn_hp'
+WK2 = '-1.39571e-08*dk2factorn_hp'
+PK2 = '1.1221778e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.01810332
+LCDSCB = -2.1685735e-09
+WCDSCB = -2.7808991e-09
+PCDSCB = 2.5748436e-16
+CDSCD = -0.034123408
+LCDSCD = 1.8392377e-09
+WCDSCD = -6.3869483e-10
+PCDSCD = 8.2621775e-17
+CIT = 0
+VOFF = -0.29344806
+LVOFF = 1.1917528e-08
+WVOFF = 1.644492e-08
+PVOFF = -1.161502e-15
+NFACTOR = 2.3640108
+LNFACTOR = -8.4270915e-08
+WNFACTOR = -1.139495e-07
+PNFACTOR = 1.0119255e-14
+ETA0 = 0
+ETAB = -0.19803551
+LETAB = 6.7296613e-09
+WETAB = -2.3369422e-09
+PETAB = 3.0230781e-16
+U0 = '(0.18072693*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.1544367e-08*du0factorn_hp'
+WU0 = '-8.3599511e-09*du0factorn_hp'
+PU0 = '7.2355829e-16*du0factorn_hp'
+UA = 4.7610771e-26
+LUA = -2.9790161e-33
+WUA = -2.5581439e-33
+PUA = 1.6050823e-40
+UB = 1e-19
+UC = -4.6916827e-27
+LUC = 2.367099e-34
+WUC = -8.2200009e-35
+PUC = 1.0633421e-41
+EU = 2.9
+VSAT = '-244193.84*dvsatfactorn_hp'
+LVSAT = '0.021246659*dvsatfactorn_hp'
+WVSAT = '0.039475574*dvsatfactorn_hp'
+PVSAT = '-2.1213717e-09*dvsatfactorn_hp'
+A0 = 4.445995
+LA0 = -2.2346745e-07
+WA0 = 7.7601344e-08
+PA0 = -1.003854e-14
+AGS = -13.82601
+LAGS = 1.235277e-06
+WAGS = 1.0378207e-06
+PAGS = -8.6469387e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.018246779
+LKETA = -3.6784728e-09
+WKETA = 1.2773927e-09
+PKETA = -1.6524377e-16
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = -0.22478226
+LPDIBLC2 = 1.7994969e-08
+WPDIBLC2 = 2.0306859e-08
+PPDIBLC2 = -1.3672475e-15
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.54123352
+LPVAG = -1.8392338e-08
+WPVAG = 6.38699e-09
+PPVAG = -8.262207e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.835645
+LPDITSD = 8.8590128e-09
+WPDITSD = -3.0747343e-09
+PPDITSD = 3.9781762e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -3.2370259e-10
+LALPHA0 = 5.5177158e-17
+WALPHA0 = -1.9160814e-17
+PALPHA0 = 2.478651e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.00975279
+LAIGC = 3.8594475e-11
+WAIGC = 4.5495353e-11
+PAIGC = -4.1811444e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 143093.35
+LAT = -0.0084547374
+WAT = -0.0088438678
+PAT = 8.0320005e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.008 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.365+dvth0n008_hp+(mcm_NENHHP_vth0*mcmScale)'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011903287
+LCDSCB = 6.5456963e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.105
+NFACTOR = -0.22582131
+LNFACTOR = 1.6364238e-07
+ETA0 = -0.34171267
+LETA0 = 3.2401196e-08
+ETAB = -0.0731796
+U0 = '(0.036403287*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.5456963e-10*du0factorn_hp'
+UA = 3.7719339e-27
+LUA = -2.6169693e-34
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '66935.181*dvsatfactorn_hp'
+LVSAT = '0.0029455655*dvsatfactorn_hp'
+A0 = 1.2216104
+LA0 = 2.7819206e-08
+AGS = 1.6903287
+LAGS = -6.5456963e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.099032866
+LKETA = -6.5456963e-09
+DWG = 0
+DWB = 0
+PCLM = 4.2341346
+LPCLM = -2.5925065e-07
+PDIBLC1 = 0
+PDIBLC2 = -0.038165073
+LPDIBLC2 = 5.9893122e-09
+PDIBLCB = -0.28554856
+LPDIBLCB = 3.6557714e-08
+DROUT = 0.56
+PVAG = 2.6363718
+LPVAG = -1.8360678e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.3549298e-10
+LALPHA0 = 9.8185444e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010095487
+LAIGC = 3.2726106e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+LVTH0 = '0.0+dlvth0n008_hp'
+WVTH0 = '0.0+dwvth0n008_hp'
+PVTH0 = '0.0+dpvth0n008_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.108 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.38607348+dvth0n108_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-2.7124469e-09+dlvth0n108_hp'
+WVTH0 = '-2.0921755e-07+dwvth0n108_hp'
+PVTH0 = '2.6929173e-14+dpvth0n108_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12826757*dk2factorn_hp'
+LK2 = '-3.4076052e-10*dk2factorn_hp'
+WK2 = '-6.6839517e-08*dk2factorn_hp'
+PK2 = '3.3830705e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.011610116
+LCDSCB = -9.7975525e-10
+WCDSCB = -2.3344106e-07
+PCDSCB = 1.6225577e-14
+CDSCD = 0.0185599
+LCDSCD = -1.363039e-09
+WCDSCD = -1.8426269e-07
+PCDSCD = 1.3532252e-14
+CIT = 0
+VOFF = -0.11006111
+LVOFF = 1.6010392e-09
+WVOFF = 5.0246707e-08
+PVOFF = -1.5895117e-14
+NFACTOR = -0.72375701
+LNFACTOR = 2.0707746e-07
+WNFACTOR = 4.9435056e-06
+PNFACTOR = -4.3122349e-13
+ETA0 = -0.34240279
+LETA0 = 3.2466632e-08
+WETA0 = 6.8514375e-09
+PETA0 = -6.4965362e-16
+ETAB = -0.0731796
+U0 = '(0.035880513*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.2404348e-10*du0factorn_hp'
+WU0 = '5.1900935e-09*du0factorn_hp'
+PU0 = '6.8973642e-16*du0factorn_hp'
+UA = 2.8495127e-27
+LUA = -1.9407349e-34
+WUA = 9.1577972e-33
+PUA = -6.7136551e-40
+UB = 1e-19
+UC = 4.6364352e-28
+LUC = -4.0891173e-35
+WUC = -6.7743064e-33
+PUC = 4.0596756e-40
+EU = 2.9
+VSAT = '69328.962*dvsatfactorn_hp'
+LVSAT = '0.002678906*dvsatfactorn_hp'
+WVSAT = '-0.023765458*dvsatfactorn_hp'
+PVSAT = '2.647395e-09*dvsatfactorn_hp'
+A0 = 1.0988302
+LA0 = 3.9461219e-08
+WA0 = 1.2189613e-06
+PA0 = -1.1558191e-13
+AGS = 1.9792232
+LAGS = -9.2849939e-08
+WAGS = -2.8681446e-06
+PAGS = 2.7195747e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.12792232
+LKETA = -9.2849939e-09
+WKETA = -2.8681446e-07
+PKETA = 2.7195747e-14
+DWG = 0
+DWB = 0
+PCLM = 4.2396562
+LPCLM = -2.5977421e-07
+WPCLM = -5.4818116e-08
+PPCLM = 5.1979029e-15
+PDIBLC1 = 0
+PDIBLC2 = -0.038292641
+LPDIBLC2 = 6.0014081e-09
+WPDIBLC2 = 1.2664951e-09
+PPDIBLC2 = -1.2008888e-16
+PDIBLCB = -0.28632722
+LPDIBLCB = 3.6631546e-08
+WPDIBLCB = 7.7305057e-09
+PPDIBLCB = -7.3300359e-16
+DROUT = 0.56
+PVAG = 3.0114805
+LPVAG = -2.1123836e-07
+WPVAG = -3.7240786e-06
+PPVAG = 2.7432641e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.3758423e-10
+LALPHA0 = 9.8383737e-17
+WALPHA0 = 2.0761947e-17
+PALPHA0 = -1.9686473e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010003164
+LAIGC = 1.2820292e-11
+WAIGC = 9.1657779e-10
+PAIGC = -9.4789382e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.208 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26164328+dvth0n208_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.0820319e-08+dlvth0n208_hp'
+WVTH0 = '1.5523852e-07+dwvth0n208_hp'
+PVTH0 = '-1.2708297e-14+dpvth0n208_hp'
+K1 = '0.59842774*dk1factorn_hp'
+LK1 = '4.9725775e-09*dk1factorn_hp'
+WK1 = '1.5691316e-07*dk1factorn_hp'
+PK1 = '-1.456468e-14*dk1factorn_hp'
+K2 = '-0.11925873*dk2factorn_hp'
+LK2 = '-1.8082179e-09*dk2factorn_hp'
+WK2 = '-9.3226432e-08*dk2factorn_hp'
+PK2 = '7.6812533e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.083339224
+LCDSCB = 5.6272004e-09
+WCDSCB = 4.4665555e-08
+PCDSCB = -3.1261957e-15
+CDSCD = -0.04595956
+LCDSCD = 3.4384275e-09
+WCDSCD = 4.7148136e-09
+PCDSCD = -5.3124381e-16
+CIT = 0
+VOFF = -0.025764541
+LVOFF = -8.9404252e-09
+WVOFF = -1.9665795e-07
+PVOFF = 1.4980832e-14
+NFACTOR = 0.6459818
+LNFACTOR = 8.5435924e-08
+WNFACTOR = 9.3154061e-07
+PNFACTOR = -7.493542e-14
+ETA0 = -0.35599965
+LETA0 = 3.4040433e-08
+WETA0 = 4.6676663e-08
+PETA0 = -5.2593143e-15
+ETAB = -0.0035737308
+LETAB = -4.8807636e-09
+WETAB = -2.0387559e-07
+PETAB = 1.4295757e-14
+U0 = '(0.027875653*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.8458407e-10*du0factorn_hp'
+WU0 = '2.8636328e-08*du0factorn_hp'
+PU0 = '-2.2645337e-15*du0factorn_hp'
+UA = 5.665269e-27
+LUA = -4.2017978e-34
+WUA = 9.1044715e-34
+PUA = -9.1001894e-42
+UB = 1e-19
+UC = 2.3893876e-27
+LUC = -1.9248482e-34
+WUC = -1.2414811e-32
+PUC = 8.4998536e-40
+EU = 2.9
+VSAT = '65151.405*dvsatfactorn_hp'
+LVSAT = '0.0033821018*dvsatfactorn_hp'
+WVSAT = '-0.011529393*dvsatfactorn_hp'
+PVSAT = '5.8773464e-10*dvsatfactorn_hp'
+A0 = 1.515
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.096788548
+LKETA = -5.3356552e-09
+WKETA = -1.9562366e-07
+PKETA = 1.5628134e-14
+DWG = 0
+DWB = 0
+PCLM = 4.3484492
+LPCLM = -2.7236667e-07
+WPCLM = -3.7347277e-07
+PPCLM = 4.2081204e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.031294345
+LPDIBLC2 = 5.6253653e-09
+WPDIBLC2 = -1.9231513e-08
+PPDIBLC2 = 9.8134048e-16
+PDIBLCB = -0.11143527
+LPDIBLCB = 2.5068096e-08
+WPDIBLCB = -5.04528e-07
+PPDIBLCB = 3.3136342e-14
+DROUT = 0.56
+PVAG = 2.2662691
+LPVAG = -1.5894238e-07
+WPVAG = -1.5413545e-06
+PPVAG = 1.2115148e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.091616
+LPDITSD = -6.424123e-09
+WPDITSD = -2.6834365e-07
+PPDITSD = 1.8816256e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.7878688e-10
+LALPHA0 = 1.0315283e-16
+WALPHA0 = 1.4144448e-16
+PALPHA0 = -1.5937321e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010306729
+LAIGC = -1.929625e-11
+WAIGC = 2.74361e-11
+PAIGC = -7.2002982e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.308 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.46305282+dvth0n308_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.0100054e-09+dlvth0n308_hp'
+WVTH0 = '-3.2072354e-08+dwvth0n308_hp'
+PVTH0 = '2.013904e-15+dpvth0n308_hp'
+K1 = '0.75793836*dk1factorn_hp'
+LK1 = '-9.7240945e-09*dk1factorn_hp'
+WK1 = '8.5682864e-09*dk1factorn_hp'
+PK1 = '-8.967746e-16*dk1factorn_hp'
+K2 = '-0.16759604*dk2factorn_hp'
+LK2 = '2.9860151e-09*dk2factorn_hp'
+WK2 = '-4.8272732e-08*dk2factorn_hp'
+PK2 = '3.2226165e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.033358771
+LCDSCB = 2.0612965e-09
+WCDSCB = -1.8162664e-09
+PCDSCB = 1.9009486e-16
+CDSCD = -0.038418395
+LCDSCD = 2.6085279e-09
+WCDSCD = -2.29847e-09
+PCDSCD = 2.4056277e-16
+CIT = 0
+VOFF = -0.3081215
+LVOFF = 1.3794303e-08
+WVOFF = 6.5934028e-08
+PVOFF = -6.1624651e-15
+NFACTOR = 2.4313257
+LNFACTOR = -5.2433565e-08
+WNFACTOR = -7.2882923e-07
+PNFACTOR = 5.3283205e-14
+ETA0 = -0.57109039
+LETA0 = 5.300861e-08
+WETA0 = 2.4671105e-07
+PETA0 = -2.289972e-14
+ETAB = -0.21375289
+LETAB = 9.5446598e-09
+WETAB = -8.4089763e-09
+PETAB = 8.8011277e-16
+U0 = '(0.064141999*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.5055716e-09*du0factorn_hp'
+WU0 = '-5.0913734e-09*du0factorn_hp'
+PU0 = '3.3031109e-16*du0factorn_hp'
+UA = 5.9446552e-27
+LUA = -3.6031115e-34
+WUA = 6.5061795e-34
+PUA = -6.4778021e-41
+UB = 1e-19
+UC = -5.0260618e-27
+LUC = 2.7196561e-34
+WUC = -5.518443e-33
+PUC = 4.1804646e-40
+EU = 2.9
+VSAT = '71821.072*dvsatfactorn_hp'
+LVSAT = '0.0014552328*dvsatfactorn_hp'
+WVSAT = '-0.017732184*dvsatfactorn_hp'
+PVSAT = '2.3797228e-09*dvsatfactorn_hp'
+A0 = 1.515
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.068974781
+LKETA = 1.0434111e-08
+WKETA = -4.1463762e-08
+PKETA = 9.6225125e-16
+DWG = 0
+DWB = 0
+PCLM = 6.7565928
+LPCLM = -4.2413614e-07
+WPCLM = -2.6130464e-06
+PPCLM = 1.8322681e-13
+PDIBLC1 = 0
+PDIBLC2 = -0.15393512
+LPDIBLC2 = 1.3873585e-08
+WPDIBLC2 = 9.4824411e-08
+PPDIBLC2 = -6.6895042e-15
+PDIBLCB = -1.4049824
+LPDIBLCB = 1.1336206e-07
+WPDIBLCB = 6.9847087e-07
+PPDIBLCB = -4.8977047e-14
+DROUT = 0.56
+PVAG = 0.5841839
+LPVAG = -2.6085275e-08
+WPVAG = 2.2984746e-08
+PPVAG = -2.4056316e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.814976
+LPDITSD = 1.2562779e-08
+WPDITSD = -1.1067952e-08
+PPDITSD = 1.1584374e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -4.5255179e-10
+LALPHA0 = 7.8255832e-17
+WALPHA0 = -6.8954148e-17
+PALPHA0 = 7.2168871e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010143324
+LAIGC = -1.7844617e-12
+WAIGC = 1.7940267e-10
+PAIGC = -1.7005993e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.8821587
+LUTE = 3.0479257e-08
+WUTE = 3.916776e-07
+PUTE = -2.8345709e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.408 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.40503071+dvth0n408_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '6.6311021e-10+dlvth0n408_hp'
+WVTH0 = '-7.0068041e-09+dwvth0n408_hp'
+PVTH0 = '-4.3688195e-16+dpvth0n408_hp'
+K1 = '0.78304577*dk1factorn_hp'
+LK1 = '-1.2874777e-08*dk1factorn_hp'
+WK1 = '-2.2781181e-09*dk1factorn_hp'
+PK1 = '4.6432047e-16*dk1factorn_hp'
+K2 = '-0.32295682*dk2factorn_hp'
+LK2 = '1.4292153e-08*dk2factorn_hp'
+WK2 = '1.8843123e-08*dk2factorn_hp'
+PK2 = '-1.6616351e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.055937055
+LCDSCB = 3.8682442e-09
+WCDSCB = 7.9375522e-09
+PCDSCB = -5.9050655e-16
+CDSCD = -0.045153538
+LCDSCD = 3.4537094e-09
+WCDSCD = 6.1111156e-10
+PCDSCD = -1.245556e-16
+CIT = 0
+VOFF = -0.16521678
+LVOFF = -8.7570638e-10
+WVOFF = 4.1991896e-09
+PVOFF = 1.7497885e-16
+NFACTOR = -0.37016079
+LNFACTOR = 1.5919683e-07
+WNFACTOR = 4.8141294e-07
+PNFACTOR = -3.8141125e-14
+ETA0 = 0
+ETAB = -0.23839411
+LETAB = 1.2636917e-08
+WETAB = 2.2360323e-09
+PETAB = -4.5574224e-16
+U0 = '(0.053344685*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.8995405e-09*du0factorn_hp'
+WU0 = '-4.2693399e-10*du0factorn_hp'
+PU0 = '6.8505634e-17*du0factorn_hp'
+UA = 4.3380227e-27
+LUA = -3.2753834e-34
+WUA = 1.3446832e-33
+PUA = -7.8935874e-41
+UB = 1e-19
+UC = -2.4201658e-26
+LUC = 1.7385702e-33
+WUC = 2.7654143e-33
+PUC = -2.1552671e-40
+EU = 2.9
+VSAT = '-20639.272*dvsatfactorn_hp'
+LVSAT = '0.01087906*dvsatfactorn_hp'
+WVSAT = '0.022210685*dvsatfactorn_hp'
+PVSAT = '-1.6913707e-09*dvsatfactorn_hp'
+A0 = 1.515
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.12615574
+LKETA = 9.9549582e-09
+WKETA = -1.6761587e-08
+PKETA = 1.1692454e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.066285954
+LPDIBLC2 = -1.7581525e-09
+WPDIBLC2 = -3.1109446e-10
+PPDIBLC2 = 6.3406588e-17
+PDIBLCB = 0.21185309
+LPDIBLCB = -1.1709837e-11
+WPDIBLCB = -2.0786003e-12
+PPDIBLCB = 4.2280164e-19
+DROUT = 0.56
+PVAG = 0.65153548
+LPVAG = -3.4537102e-08
+WPVAG = -6.1111355e-09
+PPVAG = 1.2455576e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.782545
+LPDITSD = 1.6632699e-08
+WPDITSD = 2.9419801e-09
+PPDITSD = -5.997681e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.5460619e-10
+LALPHA0 = 1.0361128e-16
+WALPHA0 = 1.8333353e-17
+PALPHA0 = -3.7366686e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010573609
+LAIGC = -5.0688347e-11
+WAIGC = -6.4802771e-12
+PAIGC = 4.1204853e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.95979518
+LUTE = -3.8336218e-08
+WUTE = -6.7834458e-09
+PUTE = 1.3825759e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.508 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.44701966+dvth0n508_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.1894976e-09+dlvth0n508_hp'
+WVTH0 = '-1.4480837e-08+dwvth0n508_hp'
+PVTH0 = '6.0488224e-16+dpvth0n508_hp'
+K1 = '0.90559072*dk1factorn_hp'
+LK1 = '-2.2016746e-08*dk1factorn_hp'
+WK1 = '-2.4091118e-08*dk1factorn_hp'
+PK1 = '2.0915909e-15*dk1factorn_hp'
+K2 = '-0.30630857*dk2factorn_hp'
+LK2 = '1.3731539e-08*dk2factorn_hp'
+WK2 = '1.5879736e-08*dk2factorn_hp'
+PK2 = '-1.5618458e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011544095
+LCDSCB = 5.6109705e-10
+WCDSCB = 3.5605249e-11
+PCDSCB = -1.834346e-18
+CDSCD = -0.042720476
+LCDSCD = 2.8054855e-09
+WCDSCD = 1.7802662e-10
+PCDSCD = -9.1717591e-18
+CIT = 0
+VOFF = -0.16598517
+LVOFF = 5.836294e-10
+WVOFF = 4.3359628e-09
+PVOFF = -8.4782914e-17
+NFACTOR = 3.673405
+LNFACTOR = -1.4358547e-07
+WNFACTOR = -2.3834176e-07
+PNFACTOR = 1.5754124e-14
+ETA0 = 0
+ETAB = -0.22949159
+LETAB = 1.0265098e-08
+WETAB = 6.5138329e-10
+PETAB = -3.3558527e-17
+U0 = '(0.0031242534*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.2475181e-09*du0factorn_hp'
+WU0 = '8.5123029e-09*du0factorn_hp'
+PU0 = '-4.916708e-16*du0factorn_hp'
+UA = 1.830988e-27
+LUA = -1.7758316e-34
+WUA = 1.7909354e-33
+PUA = -1.056279e-40
+UB = 1e-19
+UC = -1.2223745e-26
+LUC = 7.3274602e-34
+WUC = 6.3334594e-34
+PUC = -3.649001e-41
+EU = 2.9
+VSAT = '27225.642*dvsatfactorn_hp'
+LVSAT = '0.0041932732*dvsatfactorn_hp'
+WVSAT = '0.01369073*dvsatfactorn_hp'
+PVSAT = '-5.0130061e-10*dvsatfactorn_hp'
+A0 = -2.7747089
+LA0 = 3.7672224e-07
+WA0 = 7.6356818e-07
+PA0 = -6.7056558e-14
+AGS = 5.4656654
+LAGS = -3.7207136e-07
+WAGS = -7.9488845e-07
+PAGS = 6.6228703e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.50877285
+LKETA = 4.1637671e-08
+WKETA = 5.1344258e-08
+PKETA = -4.4702775e-15
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = 0.15102726
+LPDIBLC2 = -7.1303521e-09
+WPDIBLC2 = -1.5395047e-08
+PPDIBLC2 = 1.0196581e-15
+PDIBLCB = 0.21196448
+LPDIBLCB = -2.0018667e-11
+WPDIBLCB = -2.1904784e-11
+PPDIBLCB = 1.9017734e-18
+DROUT = 0.56
+PVAG = 0.62720474
+LPVAG = -2.8054852e-08
+WPVAG = -1.7802635e-09
+PPVAG = 9.1717298e-17
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.794255
+LPDITSD = 1.3511504e-08
+WPDITSD = 8.5763739e-10
+PPDITSD = -4.4195453e-17
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -5.8161432e-10
+LALPHA0 = 8.4164568e-17
+WALPHA0 = 5.3407996e-18
+PALPHA0 = -2.7515287e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010886883
+LAIGC = -5.2859544e-11
+WAIGC = -6.2243125e-11
+PAIGC = 4.5069584e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.46785528
+LUTE = -6.5557481e-08
+WUTE = -9.4348748e-08
+PUTE = 6.2279606e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.608 NMOS
+LMIN = '1.15700000e-07+dlminn_hp'
+LMAX = '1.29000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.50762788+dvth0n608_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.2434272e-08+dlvth0n608_hp'
+WVTH0 = '-2.0238618e-08+dwvth0n608_hp'
+PVTH0 = '1.2931358e-15+dpvth0n608_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '0.0077634775*dk2factorn_hp'
+LK2 = '-1.4521348e-08*dk2factorn_hp'
+WK2 = '-1.3957109e-08*dk2factorn_hp'
+PK2 = '1.1221785e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.018103317
+LCDSCB = -2.1685733e-09
+WCDSCB = -2.7808988e-09
+PCDSCB = 2.5748434e-16
+CDSCD = -0.034123412
+LCDSCD = 1.839238e-09
+WCDSCD = -6.3869449e-10
+PCDSCD = 8.262175e-17
+CIT = 0
+VOFF = -0.29344764
+LVOFF = 1.1917497e-08
+WVOFF = 1.6444897e-08
+PVOFF = -1.1615004e-15
+NFACTOR = 2.3640172
+LNFACTOR = -8.4271388e-08
+WNFACTOR = -1.1394993e-07
+PNFACTOR = 1.0119286e-14
+ETA0 = 0
+ETAB = -0.19803565
+LETAB = 6.7296719e-09
+WETAB = -2.3369307e-09
+PETAB = 3.0230697e-16
+U0 = '(0.18072695*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.1544369e-08*du0factorn_hp'
+WU0 = '-8.3599533e-09*du0factorn_hp'
+PU0 = '7.2355846e-16*du0factorn_hp'
+UA = 4.7610764e-26
+LUA = -2.9790156e-33
+WUA = -2.5581433e-33
+PUA = 1.6050819e-40
+UB = 1e-19
+UC = -4.6916829e-27
+LUC = 2.3670992e-34
+WUC = -8.2199986e-35
+PUC = 1.063342e-41
+EU = 2.9
+VSAT = '-244193.23*dvsatfactorn_hp'
+LVSAT = '0.021246613*dvsatfactorn_hp'
+WVSAT = '0.039475523*dvsatfactorn_hp'
+PVSAT = '-2.1213679e-09*dvsatfactorn_hp'
+A0 = 4.4459926
+LA0 = -2.2346728e-07
+WA0 = 7.7601534e-08
+PA0 = -1.0038554e-14
+AGS = -13.826009
+LAGS = 1.2352769e-06
+WAGS = 1.0378206e-06
+PAGS = -8.6469385e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.01824684
+LKETA = -3.6784773e-09
+WKETA = 1.2773876e-09
+PKETA = -1.652434e-16
+DWG = 0
+DWB = 0
+PCLM = 0.7078744
+PDIBLC1 = 0
+PDIBLC2 = -0.22478229
+LPDIBLC2 = 1.7994972e-08
+WPDIBLC2 = 2.0306861e-08
+PPDIBLC2 = -1.3672476e-15
+PDIBLCB = 0.2117339
+DROUT = 0.56
+PVAG = 0.54123409
+LPVAG = -1.839238e-08
+WPVAG = 6.3869482e-09
+PPVAG = -8.2621763e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.835663
+LPDITSD = 8.8576932e-09
+WPDITSD = -3.0760808e-09
+PPDITSD = 3.9791662e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -3.2370233e-10
+LALPHA0 = 5.5177139e-17
+WALPHA0 = -1.9160839e-17
+PALPHA0 = 2.4786529e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0097527787
+LAIGC = 3.8595304e-11
+WAIGC = 4.5496819e-11
+PAIGC = -4.1812522e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 143093.34
+LAT = -0.0084547368
+WAT = -0.008843867
+PAT = 8.0319999e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.009 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.365+dvth0n009_hp+(mcm_NENHHP_vth0*mcmScale)'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011903285
+LCDSCB = 6.5456949e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.105
+NFACTOR = -0.22582346
+LNFACTOR = 1.6364257e-07
+ETA0 = -0.34171268
+LETA0 = 3.2401196e-08
+ETAB = -0.0731796
+U0 = '(0.036403276*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.545687e-10*du0factorn_hp'
+UA = 3.7719338e-27
+LUA = -2.6169692e-34
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '66935.322*dvsatfactorn_hp'
+LVSAT = '0.0029455532*dvsatfactorn_hp'
+A0 = 1.22161
+LA0 = 2.7819239e-08
+AGS = 1.6903285
+LAGS = -6.5456949e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.09903285
+LKETA = -6.5456949e-09
+DWG = 0
+DWB = 0
+PCLM = 4.2341371
+LPCLM = -2.5925086e-07
+PDIBLC1 = 0
+PDIBLC2 = -0.038165072
+LPDIBLC2 = 5.9893121e-09
+PDIBLCB = -0.28554843
+LPDIBLCB = 3.6557703e-08
+DROUT = 0.56
+PVAG = 2.6363719
+LPVAG = -1.8360678e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.3549297e-10
+LALPHA0 = 9.8185443e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010095468
+LAIGC = 3.2742431e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+LVTH0 = '0.0+dlvth0n009_hp'
+WVTH0 = '0.0+dwvth0n009_hp'
+PVTH0 = '0.0+dpvth0n009_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.109 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.38607352+dvth0n109_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-2.7124501e-09+dlvth0n109_hp'
+WVTH0 = '-2.0921791e-07+dwvth0n109_hp'
+PVTH0 = '2.6929205e-14+dpvth0n109_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12826758*dk2factorn_hp'
+LK2 = '-3.4075977e-10*dk2factorn_hp'
+WK2 = '-6.6839431e-08*dk2factorn_hp'
+PK2 = '3.383063e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.01161012
+LCDSCB = -9.7975553e-10
+WCDSCB = -2.3344108e-07
+PCDSCB = 1.6225579e-14
+CDSCD = 0.0185599
+LCDSCD = -1.3630391e-09
+WCDSCD = -1.8426269e-07
+PCDSCD = 1.3532252e-14
+CIT = 0
+VOFF = -0.11006107
+LVOFF = 1.6010355e-09
+WVOFF = 5.0246287e-08
+PVOFF = -1.5895081e-14
+NFACTOR = -0.72376073
+LNFACTOR = 2.0707779e-07
+WNFACTOR = 4.9435212e-06
+PNFACTOR = -4.3122485e-13
+ETA0 = -0.3424028
+LETA0 = 3.2466633e-08
+WETA0 = 6.8515013e-09
+PETA0 = -6.4965916e-16
+ETAB = -0.0731796
+U0 = '(0.035880499*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.2404222e-10*du0factorn_hp'
+WU0 = '5.1901321e-09*du0factorn_hp'
+PU0 = '6.8973306e-16*du0factorn_hp'
+UA = 2.8495127e-27
+LUA = -1.9407349e-34
+WUA = 9.157797e-33
+PUA = -6.7136549e-40
+UB = 1e-19
+UC = 4.6364352e-28
+LUC = -4.0891173e-35
+WUC = -6.7743065e-33
+PUC = 4.0596756e-40
+EU = 2.9
+VSAT = '69329.166*dvsatfactorn_hp'
+LVSAT = '0.0026788883*dvsatfactorn_hp'
+WVSAT = '-0.023766084*dvsatfactorn_hp'
+PVSAT = '2.6474493e-09*dvsatfactorn_hp'
+A0 = 1.0988297
+LA0 = 3.9461266e-08
+WA0 = 1.2189629e-06
+PA0 = -1.1558205e-13
+AGS = 1.9792229
+LAGS = -9.284992e-08
+WAGS = -2.868144e-06
+PAGS = 2.7195742e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.12792229
+LKETA = -9.284992e-09
+WKETA = -2.868144e-07
+PKETA = 2.7195742e-14
+DWG = 0
+DWB = 0
+PCLM = 4.2396599
+LPCLM = -2.5977454e-07
+WPCLM = -5.483124e-08
+PPCLM = 5.1990423e-15
+PDIBLC1 = 0
+PDIBLC2 = -0.038292642
+LPDIBLC2 = 6.0014083e-09
+WPDIBLC2 = 1.2665157e-09
+PPDIBLC2 = -1.2009067e-16
+PDIBLCB = -0.286327
+LPDIBLCB = 3.6631527e-08
+WPDIBLCB = 7.7296279e-09
+PPDIBLCB = -7.3292737e-16
+DROUT = 0.56
+PVAG = 3.0114805
+LPVAG = -2.1123837e-07
+WPVAG = -3.7240784e-06
+PPVAG = 2.7432639e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.3758422e-10
+LALPHA0 = 9.8383735e-17
+WALPHA0 = 2.0761883e-17
+PALPHA0 = -1.9686418e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010003133
+LAIGC = 1.2822974e-11
+WAIGC = 9.1669782e-10
+PAIGC = -9.4799803e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.209 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26164308+dvth0n209_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.0820336e-08+dlvth0n209_hp'
+WVTH0 = '1.5523885e-07+dwvth0n209_hp'
+PVTH0 = '-1.2708326e-14+dpvth0n209_hp'
+K1 = '0.59842776*dk1factorn_hp'
+LK1 = '4.9725753e-09*dk1factorn_hp'
+WK1 = '1.5691309e-07*dk1factorn_hp'
+PK1 = '-1.4564673e-14*dk1factorn_hp'
+K2 = '-0.11925874*dk2factorn_hp'
+LK2 = '-1.8082165e-09*dk2factorn_hp'
+WK2 = '-9.3226322e-08*dk2factorn_hp'
+PK2 = '7.6812437e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.083339226
+LCDSCB = 5.6272006e-09
+WCDSCB = 4.4665553e-08
+PCDSCB = -3.1261956e-15
+CDSCD = -0.045959563
+LCDSCD = 3.4384277e-09
+WCDSCD = 4.7148165e-09
+PCDSCD = -5.3124405e-16
+CIT = 0
+VOFF = -0.02576472
+LVOFF = -8.9404096e-09
+WVOFF = -1.9665772e-07
+PVOFF = 1.4980812e-14
+NFACTOR = 0.64598367
+LNFACTOR = 8.5435761e-08
+WNFACTOR = 9.3153985e-07
+PNFACTOR = -7.4935353e-14
+ETA0 = -0.35599964
+LETA0 = 3.4040431e-08
+WETA0 = 4.6676654e-08
+PETA0 = -5.2593135e-15
+ETAB = -0.0035738142
+LETAB = -4.8807564e-09
+WETAB = -2.0387535e-07
+PETAB = 1.4295735e-14
+U0 = '(0.027875658*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.8458365e-10*du0factorn_hp'
+WU0 = '2.863631e-08*du0factorn_hp'
+PU0 = '-2.2645321e-15*du0factorn_hp'
+UA = 5.665268e-27
+LUA = -4.2017969e-34
+WUA = 9.104498e-34
+PUA = -9.1004192e-42
+UB = 1e-19
+UC = 2.3893879e-27
+LUC = -1.9248485e-34
+WUC = -1.2414812e-32
+PUC = 8.4998544e-40
+EU = 2.9
+VSAT = '65151.4*dvsatfactorn_hp'
+LVSAT = '0.0033821022*dvsatfactorn_hp'
+WVSAT = '-0.011529406*dvsatfactorn_hp'
+PVSAT = '5.8773574e-10*dvsatfactorn_hp'
+A0 = 1.515
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.09678855
+LKETA = -5.3356554e-09
+WKETA = -1.9562366e-07
+PKETA = 1.5628135e-14
+DWG = 0
+DWB = 0
+PCLM = 4.3484477
+LPCLM = -2.7236654e-07
+WPCLM = -3.7347054e-07
+PPCLM = 4.2081011e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.03129434
+LPDIBLC2 = 5.6253648e-09
+WPDIBLC2 = -1.9231513e-08
+PPDIBLC2 = 9.8134049e-16
+PDIBLCB = -0.11143539
+LPDIBLCB = 2.5068106e-08
+WPDIBLCB = -5.0452788e-07
+PPDIBLCB = 3.3136332e-14
+DROUT = 0.56
+PVAG = 2.2662693
+LPVAG = -1.589424e-07
+WPVAG = -1.5413548e-06
+PPVAG = 1.2115151e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.091617
+LPDITSD = -6.4242078e-09
+WPDITSD = -2.6834651e-07
+PPDITSD = 1.8816505e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.787869e-10
+LALPHA0 = 1.0315283e-16
+WALPHA0 = 1.4144453e-16
+PALPHA0 = -1.5937324e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.01030675
+LAIGC = -1.9298091e-11
+WAIGC = 2.740354e-11
+PAIGC = -7.1720296e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.309 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.463053+dvth0n309_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.0100213e-09+dlvth0n309_hp'
+WVTH0 = '-3.207238e-08+dwvth0n309_hp'
+PVTH0 = '2.0139063e-15+dpvth0n309_hp'
+K1 = '0.75793837*dk1factorn_hp'
+LK1 = '-9.7240954e-09*dk1factorn_hp'
+WK1 = '8.5682254e-09*dk1factorn_hp'
+PK1 = '-8.9676931e-16*dk1factorn_hp'
+K2 = '-0.16759579*dk2factorn_hp'
+LK2 = '2.9859934e-09*dk2factorn_hp'
+WK2 = '-4.827287e-08*dk2factorn_hp'
+PK2 = '3.2226285e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.033358786
+LCDSCB = 2.0612978e-09
+WCDSCB = -1.8162558e-09
+PCDSCB = 1.9009394e-16
+CDSCD = -0.038418393
+LCDSCD = 2.6085278e-09
+WCDSCD = -2.298471e-09
+PCDSCD = 2.4056286e-16
+CIT = 0
+VOFF = -0.3081213
+LVOFF = 1.3794285e-08
+WVOFF = 6.5933903e-08
+PVOFF = -6.1624543e-15
+NFACTOR = 2.4313276
+LNFACTOR = -5.2433725e-08
+WNFACTOR = -7.2882996e-07
+PNFACTOR = 5.3283268e-14
+ETA0 = -0.57109038
+LETA0 = 5.3008609e-08
+WETA0 = 2.4671105e-07
+PETA0 = -2.2899719e-14
+ETAB = -0.21375247
+LETAB = 9.544624e-09
+WETAB = -8.4091932e-09
+PETAB = 8.801316e-16
+U0 = '(0.064141968*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.5055689e-09*du0factorn_hp'
+WU0 = '-5.0913581e-09*du0factorn_hp'
+PU0 = '3.3030976e-16*du0factorn_hp'
+UA = 5.9446599e-27
+LUA = -3.6031155e-34
+WUA = 6.5061526e-34
+PUA = -6.4777786e-41
+UB = 1e-19
+UC = -5.0260635e-27
+LUC = 2.7196576e-34
+WUC = -5.518442e-33
+PUC = 4.1804637e-40
+EU = 2.9
+VSAT = '71821.012*dvsatfactorn_hp'
+LVSAT = '0.001455238*dvsatfactorn_hp'
+WVSAT = '-0.017732145*dvsatfactorn_hp'
+PVSAT = '2.3797194e-09*dvsatfactorn_hp'
+A0 = 1.515
+AGS = 1
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.068974782
+LKETA = 1.0434111e-08
+WKETA = -4.1463764e-08
+PKETA = 9.6225144e-16
+DWG = 0
+DWB = 0
+PCLM = 6.7565945
+LPCLM = -4.2413628e-07
+WPCLM = -2.6130471e-06
+PPCLM = 1.8322687e-13
+PDIBLC1 = 0
+PDIBLC2 = -0.1539351
+LPDIBLC2 = 1.3873584e-08
+WPDIBLC2 = 9.4824398e-08
+PPDIBLC2 = -6.689503e-15
+PDIBLCB = -1.4049824
+LPDIBLCB = 1.1336206e-07
+WPDIBLCB = 6.984708e-07
+PPDIBLCB = -4.8977041e-14
+DROUT = 0.56
+PVAG = 0.58418378
+LPVAG = -2.6085264e-08
+WPVAG = 2.2984711e-08
+PPVAG = -2.4056286e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.814985
+LPDITSD = 1.2562004e-08
+WPDITSD = -1.1078205e-08
+PPDITSD = 1.1593276e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -4.5255178e-10
+LALPHA0 = 7.8255831e-17
+WALPHA0 = -6.8954133e-17
+PALPHA0 = 7.2168858e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010143302
+LAIGC = -1.7825545e-12
+WAIGC = 1.7941026e-10
+PAIGC = -1.7006652e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.8821578
+LUTE = 3.0479182e-08
+WUTE = 3.9167678e-07
+PUTE = -2.8345639e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.409 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.49044216+dvth0n409_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.7523118e-09+dlvth0n409_hp'
+WVTH0 = '-4.3904497e-08+dwvth0n409_hp'
+PVTH0 = '2.7665758e-15+dpvth0n409_hp'
+K1 = '0.86591181*dk1factorn_hp'
+LK1 = '-2.0069207e-08*dk1factorn_hp'
+WK1 = '-3.8076302e-08*dk1factorn_hp'
+PK1 = '3.5723188e-15*dk1factorn_hp'
+K2 = '-0.36296949*dk2factorn_hp'
+LK2 = '1.7766054e-08*dk2factorn_hp'
+WK2 = '3.612857e-08*dk2factorn_hp'
+PK2 = '-3.1623576e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.06038288
+LCDSCB = 4.2542308e-09
+WCDSCB = 9.8581526e-09
+PCDSCB = -7.5725307e-16
+CDSCD = -0.083471567
+LCDSCD = 6.7804807e-09
+WCDSCD = 1.71645e-08
+PCDSCD = -1.5617208e-15
+CIT = 0
+VOFF = -0.20933653
+LVOFF = 2.9547697e-09
+WVOFF = 2.3258881e-08
+PVOFF = -1.4797836e-15
+NFACTOR = 0.87886447
+LNFACTOR = 5.0756454e-08
+WNFACTOR = -5.816591e-08
+PNFACTOR = 8.7051113e-15
+ETA0 = 0
+ETAB = -0.37859753
+LETAB = 2.4809378e-08
+WETAB = 6.2803871e-08
+PETAB = -5.714242e-15
+U0 = '(0.070397408*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.3800579e-09*du0factorn_hp'
+WU0 = '-7.7937085e-09*du0factorn_hp'
+PU0 = '7.08089e-16*du0factorn_hp'
+UA = 1.2173408e-26
+LUA = -1.0078065e-33
+WUA = -2.0402039e-33
+PUA = 2.1494002e-40
+UB = 1e-19
+UC = -3.1658327e-26
+LUC = 2.3859582e-33
+WUC = 5.9866958e-33
+PUC = -4.9519837e-40
+EU = 2.9
+VSAT = '423.7683*dvsatfactorn_hp'
+LVSAT = '0.0090503673*dvsatfactorn_hp'
+WVSAT = '0.013111464*dvsatfactorn_hp'
+PVSAT = '-9.0137638e-10*dvsatfactorn_hp'
+A0 = 1.7000207
+LA0 = -1.6063496e-08
+WA0 = -7.9928936e-08
+PA0 = 6.9394302e-15
+AGS = 1.6435529
+LAGS = -5.587326e-08
+WAGS = -2.7801484e-07
+PAGS = 2.4137248e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.35606393
+LKETA = 2.9915587e-08
+WKETA = 8.2558748e-08
+PKETA = -7.4537461e-15
+DWG = 0
+DWB = 0
+PCLM = -0.98131153
+LPCLM = 1.4665512e-07
+WPCLM = 7.2972832e-07
+PPCLM = -6.3355013e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.13534577
+LPDIBLC2 = -7.7539257e-09
+WPDIBLC2 = -3.014494e-08
+PPDIBLC2 = 2.653581e-15
+PDIBLCB = 0.39169504
+LPDIBLCB = -1.5625588e-08
+WPDIBLCB = -7.7693837e-08
+PPDIBLCB = 6.7456213e-15
+DROUT = 0.56
+PVAG = 0.39116253
+LPVAG = -1.1931522e-08
+WPVAG = 1.0636989e-07
+PPVAG = -8.5200451e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.597975
+LPDITSD = 3.2657124e-08
+WPDITSD = 8.2670109e-08
+PPDITSD = -7.5217642e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -9.9970586e-10
+LALPHA0 = 1.3357284e-16
+WALPHA0 = 1.6741643e-16
+PALPHA0 = -1.6680061e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.015173347
+LAIGBINV = 4.1905e-10
+WAIGBINV = 2.085114e-09
+PAIGBINV = -1.810296e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010795893
+LAIGC = -6.9987068e-11
+WAIGC = -1.0250899e-10
+PAIGC = 1.2457698e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.71305275
+LUTE = -5.9758395e-08
+WUTE = -1.1337661e-07
+PUTE = 1.0636994e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.509 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.23760479+dvth0n509_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.2991901e-08+dlvth0n509_hp'
+WVTH0 = '1.1005542e-09+dwvth0n509_hp'
+PVTH0 = '-7.4789413e-16+dpvth0n509_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14746253*dk2factorn_hp'
+LK2 = '-5.9474693e-11*dk2factorn_hp'
+WK2 = '-2.2316705e-09*dk2factorn_hp'
+PK2 = '1.0586495e-17*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0032346885
+LCDSCB = -1.6032559e-10
+WCDSCB = -3.1422544e-10
+PCDSCB = 2.8537954e-17
+CDSCD = 0.028226013
+LCDSCD = -3.3540887e-09
+WCDSCD = -2.7176691e-09
+PCDSCD = 2.4223255e-16
+CIT = 0
+VOFF = -0.055442881
+LVOFF = -9.0136523e-09
+WVOFF = -4.1341877e-09
+PVOFF = 6.5059556e-16
+NFACTOR = 0.065801177
+LNFACTOR = 1.6962669e-07
+WNFACTOR = 8.6559356e-08
+PNFACTOR = -1.2453791e-14
+ETA0 = 0
+ETAB = 0.030096893
+LETAB = -1.2272374e-08
+WETAB = -9.9437361e-09
+PETAB = 8.8630974e-16
+U0 = '(0.008773879*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '7.5701765e-10*du0factorn_hp'
+WU0 = '3.1752797e-09*du0factorn_hp'
+PU0 = '-2.8310441e-17*du0factorn_hp'
+UA = -2.2232884e-27
+LUA = 1.7440911e-34
+WUA = 5.2240808e-34
+PUA = 4.5056461e-42
+UB = 1e-19
+UC = 5.2296945e-27
+LUC = -7.8256162e-34
+WUC = -5.7937201e-34
+PUC = 6.8798163e-41
+EU = 2.9
+VSAT = '11048.451*dvsatfactorn_hp'
+LVSAT = '0.005597777*dvsatfactorn_hp'
+WVSAT = '0.01122027*dvsatfactorn_hp'
+PVSAT = '-2.8681531e-10*dvsatfactorn_hp'
+A0 = 0.10448089
+LA0 = 1.2675098e-07
+WA0 = 2.0407715e-07
+PA0 = -1.8481547e-14
+AGS = 0.7154008
+LAGS = 4.034661e-08
+WAGS = -1.1280377e-07
+PAGS = 7.0101113e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.18825228
+LKETA = -1.8878051e-08
+WKETA = -1.4329538e-08
+PKETA = 1.2315215e-15
+DWG = 0
+DWB = 0
+PCLM = 3.7945601
+LPCLM = -2.6798605e-07
+WPCLM = -1.2037682e-07
+PPCLM = 1.0451116e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.060817075
+LPDIBLC2 = 1.1261973e-08
+WPDIBLC2 = 4.7720468e-09
+PPDIBLC2 = -7.3124891e-16
+PDIBLCB = -0.11675791
+LPDIBLCB = 2.8519659e-08
+WPDIBLCB = 1.2810788e-08
+PPDIBLCB = -1.1122326e-15
+DROUT = 0.56
+PVAG = 1.0937176
+LPVAG = -6.8557503e-08
+WPVAG = -1.8684919e-08
+PPVAG = 1.5593795e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.135949
+LPDITSD = -1.6154378e-08
+WPDITSD = -1.3089364e-08
+PPDITSD = 1.1666832e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 7.6808037e-11
+LALPHA0 = 2.7000339e-17
+WALPHA0 = -2.4203044e-17
+PALPHA0 = 2.2898437e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.028819861
+LAIGBINV = -7.657403e-10
+WAIGBINV = -3.4396537e-10
+PAIGBINV = 2.9863073e-17
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010160397
+LAIGC = 1.0214034e-11
+WAIGC = 1.0609402e-11
+PAIGC = -1.818098e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4431348
+LUTE = 1.9116285e-08
+WUTE = 1.657799e-08
+PUTE = -3.4026988e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.609 NMOS
+LMIN = '1.29000000e-07+dlminn_hp'
+LMAX = '1.33000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.335107+dvth0n609_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.5439903e-09+dlvth0n609_hp'
+WVTH0 = '-8.1621557e-09+dwvth0n609_hp'
+PVTH0 = '2.446574e-16+dpvth0n609_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11307761*dk2factorn_hp'
+LK2 = '-4.029925e-09*dk2factorn_hp'
+WK2 = '-5.4982375e-09*dk2factorn_hp'
+PK2 = '3.8777927e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.035685833
+LCDSCB = -3.6950873e-09
+WCDSCB = -4.011675e-09
+PCDSCB = 3.6434032e-16
+CDSCD = 0.11964542
+LCDSCD = -1.1510972e-08
+WCDSCD = -1.1402512e-08
+PCDSCD = 1.0171364e-15
+CIT = 0
+VOFF = -0.21219302
+LVOFF = 4.8629705e-09
+WVOFF = 1.0757075e-08
+PVOFF = -6.6768361e-16
+NFACTOR = 1.6511672
+LNFACTOR = -2.2381748e-08
+WNFACTOR = -6.4050415e-08
+PNFACTOR = 5.7870108e-15
+ETA0 = 0
+ETAB = 0.36459612
+LETAB = -4.2118018e-08
+WETAB = -4.1721162e-08
+PETAB = 3.721646e-15
+U0 = '(-0.011285395*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '5.1261432e-09*du0factorn_hp'
+WU0 = '5.0809108e-09*du0factorn_hp'
+PU0 = '-4.4337736e-16*du0factorn_hp'
+UA = -1.8536577e-26
+LUA = 2.7638965e-33
+WUA = 2.0721705e-33
+PUA = -2.4149566e-40
+UB = 1e-19
+UC = 1.3122672e-26
+LUC = -1.3099324e-33
+WUC = -1.3292049e-33
+PUC = 1.1889839e-40
+EU = 2.9
+VSAT = '-404485.3*dvsatfactorn_hp'
+LVSAT = '0.035163171*dvsatfactorn_hp'
+WVSAT = '0.050695977*dvsatfactorn_hp'
+PVSAT = '-3.0955277e-09*dvsatfactorn_hp'
+A0 = -6.9927243
+LA0 = 7.6964212e-07
+WA0 = 8.7831164e-07
+PA0 = -7.9556205e-14
+AGS = -4.5936278
+LAGS = 4.3372157e-07
+WAGS = 3.9155395e-07
+PAGS = -3.036051e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.039990476
+LKETA = -5.5662598e-09
+WKETA = -2.4466634e-10
+PKETA = -3.3098671e-17
+DWG = 0
+DWB = 0
+PCLM = 7.622207
+LPCLM = -6.0030236e-07
+WPCLM = -4.8400328e-07
+PPCLM = 4.2021165e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.22310704
+LPDIBLC2 = 1.7849526e-08
+WPDIBLC2 = 2.0189593e-08
+PPDIBLC2 = -1.3570665e-15
+PDIBLCB = -0.52410345
+LPDIBLCB = 6.3885399e-08
+WPDIBLCB = 5.1508615e-08
+PPDIBLCB = -4.4719779e-15
+DROUT = 0.56
+PVAG = 1.6377972
+LPVAG = -1.1359599e-07
+WPVAG = -7.0372475e-08
+PPVAG = 5.8380355e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.57621
+LPDITSD = -5.5436622e-08
+WPDITSD = -5.4914133e-08
+PPDITSD = 4.8984963e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 9.9654865e-10
+LALPHA0 = -5.9447051e-17
+WALPHA0 = -1.115784e-16
+PALPHA0 = 1.0502346e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.039756856
+LAIGBINV = -1.7152902e-09
+WAIGBINV = -1.3829799e-09
+PAIGBINV = 1.2007031e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0099062036
+LAIGC = 2.5274949e-11
+WAIGC = 3.4757736e-11
+PAIGC = -3.248885e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.72999254
+LUTE = -6.3466067e-08
+WUTE = -5.1170522e-08
+PUTE = 4.4426247e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 143093.31
+LAT = -0.0084547344
+WAT = -0.0088438644
+PAT = 8.0319976e-10
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.010 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.365+dvth0n010_hp+(mcm_NENHHP_vth0*mcmScale)'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.011903287
+LCDSCB = 6.545697e-10
+CDSCD = 0
+CIT = 0
+VOFF = -0.105
+NFACTOR = -0.22582067
+LNFACTOR = 1.6364232e-07
+ETA0 = -0.34171268
+LETA0 = 3.2401196e-08
+ETAB = -0.0731796
+U0 = '(0.036403296*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.5457056e-10*du0factorn_hp'
+UA = 3.771934e-27
+LUA = -2.6169694e-34
+UB = 1e-19
+UC = -2.187e-28
+EU = 2.9
+VSAT = '66935.201*dvsatfactorn_hp'
+LVSAT = '0.0029455643*dvsatfactorn_hp'
+A0 = 1.2216105
+LA0 = 2.7819189e-08
+AGS = 1.6903287
+LAGS = -6.545697e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.099032872
+LKETA = -6.545697e-09
+DWG = 0
+DWB = 0
+PCLM = 4.2341338
+LPCLM = -2.5925057e-07
+PDIBLC1 = 0
+PDIBLC2 = -0.03816506
+LPDIBLC2 = 5.989311e-09
+PDIBLCB = -0.28554861
+LPDIBLCB = 3.6557719e-08
+DROUT = 0.56
+PVAG = 2.6363719
+LPVAG = -1.8360678e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.3549286e-10
+LALPHA0 = 9.8185433e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010095488
+LAIGC = 3.2723899e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+LVTH0 = '0.0+dlvth0n010_hp'
+WVTH0 = '0.0+dwvth0n010_hp'
+PVTH0 = '0.0+dpvth0n010_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.110 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.38607345+dvth0n110_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-2.712444e-09+dlvth0n110_hp'
+WVTH0 = '-2.0921724e-07+dwvth0n110_hp'
+PVTH0 = '2.6929144e-14+dpvth0n110_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12826757*dk2factorn_hp'
+LK2 = '-3.4076056e-10*dk2factorn_hp'
+WK2 = '-6.6839517e-08*dk2factorn_hp'
+PK2 = '3.3830709e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.011610115
+LCDSCB = -9.7975515e-10
+WCDSCB = -2.3344106e-07
+PCDSCB = 1.6225577e-14
+CDSCD = 0.018559899
+LCDSCD = -1.363039e-09
+WCDSCD = -1.8426268e-07
+PCDSCD = 1.3532251e-14
+CIT = 0
+VOFF = -0.11006111
+LVOFF = 1.6010395e-09
+WVOFF = 5.0246716e-08
+PVOFF = -1.589512e-14
+NFACTOR = -0.72375591
+LNFACTOR = 2.0707735e-07
+WNFACTOR = 4.943501e-06
+PNFACTOR = -4.3122302e-13
+ETA0 = -0.34240279
+LETA0 = 3.2466633e-08
+WETA0 = 6.8514532e-09
+PETA0 = -6.4965479e-16
+ETAB = -0.0731796
+U0 = '(0.035880532*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.2404528e-10*du0factorn_hp'
+WU0 = '5.1900005e-09*du0factorn_hp'
+PU0 = '6.8974502e-16*du0factorn_hp'
+UA = 2.8495131e-27
+LUA = -1.9407353e-34
+WUA = 9.1577942e-33
+PUA = -6.7136523e-40
+UB = 1e-19
+UC = 4.6364347e-28
+LUC = -4.0891168e-35
+WUC = -6.774306e-33
+PUC = 4.0596752e-40
+EU = 2.9
+VSAT = '69328.935*dvsatfactorn_hp'
+LVSAT = '0.0026789094*dvsatfactorn_hp'
+WVSAT = '-0.02376499*dvsatfactorn_hp'
+PVSAT = '2.64735e-09*dvsatfactorn_hp'
+A0 = 1.0988305
+LA0 = 3.9461196e-08
+WA0 = 1.2189606e-06
+PA0 = -1.1558184e-13
+AGS = 1.9792233
+LAGS = -9.2849949e-08
+WAGS = -2.8681449e-06
+PAGS = 2.719575e-13
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.12792233
+LKETA = -9.2849949e-09
+WKETA = -2.8681449e-07
+PKETA = 2.719575e-14
+DWG = 0
+DWB = 0
+PCLM = 4.2396553
+LPCLM = -2.5977412e-07
+WPCLM = -5.4817286e-08
+PPCLM = 5.197775e-15
+PDIBLC1 = 0
+PDIBLC2 = -0.038292622
+LPDIBLC2 = 6.0014064e-09
+WPDIBLC2 = 1.2664293e-09
+PPDIBLC2 = -1.2008283e-16
+PDIBLCB = -0.28632728
+LPDIBLCB = 3.6631553e-08
+WPDIBLCB = 7.7306429e-09
+PPDIBLCB = -7.3301956e-16
+DROUT = 0.56
+PVAG = 3.0114805
+LPVAG = -2.1123837e-07
+WPVAG = -3.7240787e-06
+PPVAG = 2.7432642e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -6.375841e-10
+LALPHA0 = 9.8383725e-17
+WALPHA0 = 2.0761894e-17
+PALPHA0 = -1.9686428e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010003168
+LAIGC = 1.2819848e-11
+WAIGC = 9.1655867e-10
+PAIGC = -9.4787166e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.210 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29684625+dvth0n210_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '7.6231846e-09+dlvth0n210_hp'
+WVTH0 = '5.2129246e-08+dwvth0n210_hp'
+PVTH0 = '-3.3439123e-15+dpvth0n210_hp'
+K1 = '0.62521386*dk1factorn_hp'
+LK1 = '2.5398615e-09*dk1factorn_hp'
+WK1 = '7.8456595e-08*dk1factorn_hp'
+PK1 = '-7.4392543e-15*dk1factorn_hp'
+K2 = '-0.13542606*dk2factorn_hp'
+LK2 = '-3.399012e-10*dk2factorn_hp'
+WK2 = '-4.5872326e-08*dk2factorn_hp'
+PK2 = '3.3805538e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.092292263
+LCDSCB = 6.4403153e-09
+WCDSCB = 7.0889004e-08
+PCDSCB = -5.5078094e-15
+CDSCD = -0.058693813
+LCDSCD = 4.5949523e-09
+WCDSCD = 4.2013443e-08
+PCDSCD = -3.9187053e-15
+CIT = 0
+VOFF = -0.063148946
+LVOFF = -5.5451742e-09
+WVOFF = -8.7159017e-08
+PVOFF = 5.0361401e-15
+NFACTOR = 0.91123993
+LNFACTOR = 6.1345187e-08
+WNFACTOR = 1.5459819e-07
+PNFACTOR = -4.3735125e-15
+ETA0 = -0.42713598
+LETA0 = 4.0501034e-08
+WETA0 = 2.5503496e-07
+PETA0 = -2.4182414e-14
+ETAB = -0.050167885
+LETAB = -6.4908284e-10
+WETAB = -6.7401313e-08
+PETAB = 1.9011636e-15
+U0 = '(0.036316567*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.8201965e-10*du0factorn_hp'
+WU0 = '3.9128562e-09*du0factorn_hp'
+PU0 = '-1.9148052e-17*du0factorn_hp'
+UA = 6.7439136e-27
+LUA = -5.1814229e-34
+WUA = -2.2489047e-33
+PUA = 2.7783216e-40
+UB = 1e-19
+UC = -6.8288428e-28
+LUC = 8.6538915e-35
+WUC = -3.4161262e-33
+PUC = 3.2724804e-41
+EU = 2.9
+VSAT = '58421.182*dvsatfactorn_hp'
+LVSAT = '0.0039933406*dvsatfactorn_hp'
+WVSAT = '0.0081838164*dvsatfactorn_hp'
+PVSAT = '-1.2026191e-09*dvsatfactorn_hp'
+A0 = 1.5788111
+LA0 = -5.7953217e-09
+WA0 = -1.8690263e-07
+PA0 = 1.6974497e-14
+AGS = 1.2219507
+LAGS = -2.0157565e-08
+WAGS = -6.5009369e-07
+PAGS = 5.9041509e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.05694907
+LKETA = -1.7174338e-09
+WKETA = -7.8933827e-08
+PKETA = 5.0303637e-15
+DWG = 0
+DWB = 0
+PCLM = 4.7745899
+LPCLM = -3.1106877e-07
+WPCLM = -1.6216406e-06
+PPCLM = 1.5543982e-13
+PDIBLC1 = 0
+PDIBLC2 = -0.043874956
+LPDIBLC2 = 6.7679365e-09
+WPDIBLC2 = 1.7617088e-08
+PPDIBLC2 = -2.3652494e-15
+PDIBLCB = -0.31903972
+LPDIBLCB = 4.3922731e-08
+WPDIBLCB = 1.0354538e-07
+PPDIBLCB = -2.2088882e-14
+DROUT = 0.56
+PVAG = 2.171661
+LPVAG = -1.5035007e-07
+WPVAG = -1.2642473e-06
+PPVAG = 9.5984605e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.030289
+LPDITSD = -8.5435948e-10
+WPDITSD = -8.8715526e-08
+PPDITSD = 2.5024189e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -7.8337603e-10
+LALPHA0 = 1.1265162e-16
+WALPHA0 = 4.4778645e-16
+PALPHA0 = -4.3759298e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.018335371
+LAIGBINV = 1.5118156e-10
+WAIGBINV = 4.875697e-09
+PAIGBINV = -4.428108e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010301537
+LAIGC = -1.8824624e-11
+WAIGC = 4.2634804e-11
+PAIGC = -2.1005064e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4948471
+LUTE = 3.0739914e-09
+WUTE = 9.9138085e-08
+PUTE = -9.0037209e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.310 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.35019254+dvth0n310_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '5.2399662e-09+dlvth0n310_hp'
+WVTH0 = '2.5171973e-09+dwvth0n310_hp'
+PVTH0 = '-1.1275192e-15+dpvth0n310_hp'
+K1 = '0.67769325*dk1factorn_hp'
+LK1 = '-2.4362336e-09*dk1factorn_hp'
+WK1 = '2.9650769e-08*dk1factorn_hp'
+PK1 = '-2.8114859e-15*dk1factorn_hp'
+K2 = '-0.13231099*dk2factorn_hp'
+LK2 = '-2.1857235e-10*dk2factorn_hp'
+WK2 = '-4.8769341e-08*dk2factorn_hp'
+PK2 = '3.267718e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0062749919
+LCDSCB = -3.9845235e-10
+WCDSCB = -9.1070578e-09
+PCDSCB = 8.5224458e-16
+CDSCD = 0.00017527531
+LCDSCD = -8.9654922e-10
+WCDSCD = -1.273481e-08
+PCDSCD = 1.1883911e-15
+CIT = 0
+VOFF = -0.17285395
+LVOFF = 1.5093045e-09
+WVOFF = 1.4866637e-08
+PVOFF = -1.5245252e-15
+NFACTOR = 1.358823
+LNFACTOR = 4.4971135e-08
+WNFACTOR = -2.616541e-07
+PNFACTOR = 1.0854357e-14
+ETA0 = -0.28554519
+LETA0 = 2.7075395e-08
+WETA0 = 1.2335552e-07
+PETA0 = -1.1696571e-14
+ETAB = -0.072539826
+LETAB = -3.2803086e-09
+WETAB = -4.6595408e-08
+PETAB = 4.3482036e-15
+U0 = '(0.035897603*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '5.9584317e-11*du0factorn_hp'
+WU0 = '4.3024923e-09*du0factorn_hp'
+PU0 = '-5.2283974e-16*du0factorn_hp'
+UA = 2.7954316e-27
+LUA = -7.429864e-35
+WUA = 1.4231835e-33
+PUA = -1.3494243e-40
+UB = 1e-19
+UC = 2.5259624e-27
+LUC = -4.1390923e-34
+WUC = -6.4003536e-33
+PUC = 4.9814158e-40
+EU = 2.9
+VSAT = '90548.347*dvsatfactorn_hp'
+LVSAT = '-0.00024557852*dvsatfactorn_hp'
+WVSAT = '-0.021694447*dvsatfactorn_hp'
+PVSAT = '2.7395757e-09*dvsatfactorn_hp'
+A0 = 1.3187208
+LA0 = 1.7826077e-08
+WA0 = 5.498132e-08
+PA0 = -4.9934035e-15
+AGS = 0.31729605
+LAGS = 6.2003173e-08
+WAGS = 1.9123517e-07
+PAGS = -1.7367978e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.030442813
+LKETA = 1.4050055e-09
+WKETA = -5.4283008e-08
+PKETA = 2.1264951e-15
+DWG = 0
+DWB = 0
+PCLM = 4.4995082
+LPCLM = -2.191477e-07
+WPCLM = -1.3658146e-06
+PPCLM = 6.9953223e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.081028371
+LPDIBLC2 = 7.2521942e-09
+WPDIBLC2 = 5.2169763e-08
+PPDIBLC2 = -2.8156091e-15
+PDIBLCB = -0.51345916
+LPDIBLCB = 3.2393918e-08
+WPDIBLCB = 2.8435547e-07
+PPDIBLCB = -1.1367086e-14
+DROUT = 0.56
+PVAG = 0.88095097
+LPVAG = -5.303766e-08
+WPVAG = -6.3886994e-08
+PPVAG = 5.4840596e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.000838
+LPDITSD = -4.317215e-09
+WPDITSD = -6.1326466e-08
+PPDITSD = 5.7228746e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -1.4812149e-10
+LALPHA0 = 5.0607472e-17
+WALPHA0 = -1.4300027e-16
+PALPHA0 = 1.3941756e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.025120268
+LAIGBINV = -4.6502277e-10
+WAIGBINV = -1.4342571e-09
+PAIGBINV = 1.3025923e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010207227
+LAIGC = -7.5882043e-12
+WAIGC = 1.3034315e-10
+PAIGC = -1.2550377e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6650772
+LUTE = 1.0763919e-08
+WUTE = 2.5745211e-07
+PUTE = -1.6155354e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.410 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.43467006+dvth0n410_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.6870894e-09+dlvth0n410_hp'
+WVTH0 = '-3.3977092e-08+dwvth0n410_hp'
+PVTH0 = '1.8649688e-15+dpvth0n410_hp'
+K1 = '0.81243406*dk1factorn_hp'
+LK1 = '-1.5212357e-08*dk1factorn_hp'
+WK1 = '-2.8557263e-08*dk1factorn_hp'
+PK1 = '2.7077996e-15*dk1factorn_hp'
+K2 = '-0.30491215*dk2factorn_hp'
+LK2 = '1.2493286e-08*dk2factorn_hp'
+WK2 = '2.5794363e-08*dk2factorn_hp'
+PK2 = '-2.223805e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.043023048
+LCDSCB = 2.6776109e-09
+WCDSCB = 6.7681026e-09
+PCDSCB = -4.7661474e-16
+CDSCD = -0.05891989
+LCDSCD = 4.5506973e-09
+WCDSCD = 1.2794302e-08
+PCDSCD = -1.1648194e-15
+CIT = 0
+VOFF = -0.18032778
+LVOFF = 3.2019515e-10
+WVOFF = 1.8095331e-08
+PVOFF = -1.0108299e-15
+NFACTOR = 0.89403676
+LNFACTOR = 4.9378506e-08
+WNFACTOR = -6.0866427e-08
+PNFACTOR = 8.9503722e-15
+ETA0 = 0
+ETAB = -0.28876441
+LETAB = 1.6650734e-08
+WETAB = 4.6813611e-08
+PETAB = -4.2620066e-15
+U0 = '(0.059343402*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.376133e-09*du0factorn_hp'
+WU0 = '-5.826093e-09*du0factorn_hp'
+PU0 = '5.2939016e-16*du0factorn_hp'
+UA = 9.8588486e-27
+LUA = -7.9759821e-34
+WUA = -1.6282127e-33
+PUA = 1.7752298e-40
+UB = 1e-19
+UC = -2.228603e-26
+LUC = 1.5347662e-33
+WUC = 4.3184272e-33
+PUC = -3.4368621e-40
+EU = 2.9
+VSAT = '16675.575*dvsatfactorn_hp'
+LVSAT = '0.0075743782*dvsatfactorn_hp'
+WVSAT = '0.010218591*dvsatfactorn_hp'
+PVSAT = '-6.3864564e-10*dvsatfactorn_hp'
+A0 = 1.5826546
+LA0 = -5.4043119e-09
+WA0 = -5.90381e-08
+PA0 = 5.0421245e-15
+AGS = 1.2353131
+LAGS = -1.8796927e-08
+WAGS = -2.0534821e-07
+PAGS = 1.7537665e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.2374452
+LKETA = 1.9142634e-08
+WKETA = 6.1444612e-08
+PKETA = -5.5361603e-15
+DWG = 0
+DWB = 0
+PCLM = 0.090228565
+LPCLM = 4.9337851e-08
+WPCLM = 5.3899415e-07
+PPCLM = -4.6032535e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.091412983
+LPDIBLC2 = -3.76395e-09
+WPDIBLC2 = -2.2324902e-08
+PPDIBLC2 = 1.9433652e-15
+PDIBLCB = 0.27761107
+LPDIBLCB = -5.2644817e-09
+WPDIBLCB = -5.7386876e-08
+PPDIBLCB = 4.9013431e-15
+DROUT = 0.56
+PVAG = 0.5538857
+LPVAG = -2.6710041e-08
+WPVAG = 7.7405202e-08
+PPVAG = -5.889472e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.716246
+LPDITSD = 2.1915706e-08
+WPDITSD = 6.161729e-08
+PPDITSD = -5.6097472e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -7.734548e-10
+LALPHA0 = 1.1302472e-16
+WALPHA0 = 1.2714372e-16
+PALPHA0 = -1.3022493e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.018235163
+LAIGBINV = 1.4097586e-10
+WAIGBINV = 1.5401083e-09
+PAIGBINV = -1.3153218e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010711438
+LAIGC = -6.2316855e-11
+WAIGC = -8.747598e-11
+PAIGC = 1.10924e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -0.87228837
+LUTE = -4.5296616e-08
+WUTE = -8.503267e-08
+PUTE = 8.0627977e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.510 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.25492592+dvth0n510_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.1418796e-08+dlvth0n510_hp'
+WVTH0 = '-1.9826363e-09+dwvth0n510_hp'
+PVTH0 = '-4.6787877e-16+dpvth0n510_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13533024*dk2factorn_hp'
+LK2 = '-1.1613288e-09*dk2factorn_hp'
+WK2 = '-4.3912172e-09*dk2factorn_hp'
+PK2 = '2.0671653e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0.012787379
+LCDSCD = -1.9519519e-09
+WCDSCD = 3.0408072e-11
+PCDSCD = -7.3478253e-18
+CIT = 0
+VOFF = -0.063600781
+LVOFF = -8.2727519e-09
+WVOFF = -2.6820747e-09
+PVOFF = 5.1871466e-16
+NFACTOR = 0.13737458
+LNFACTOR = 1.6312639e-07
+WNFACTOR = 7.3819441e-08
+PNFACTOR = -1.1296752e-14
+ETA0 = 0
+ETAB = -0.02639152
+LETAB = -7.142096e-09
+WETAB = 1.1123713e-10
+PETAB = -2.688293e-17
+U0 = '(0.028052279*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-9.9384666e-10*du0factorn_hp'
+WU0 = '-2.5627308e-10*du0factorn_hp'
+PU0 = '2.8334318e-16*du0factorn_hp'
+UA = 4.4180047e-27
+LUA = -4.2875313e-34
+WUA = -6.5974247e-34
+PUA = 1.1186856e-40
+UB = 1e-19
+UC = 3.4411031e-27
+LUC = -6.2012175e-34
+WUC = -2.6100252e-34
+PUC = 3.9883846e-41
+EU = 2.9
+VSAT = '27141.536*dvsatfactorn_hp'
+LVSAT = '0.0041362031*dvsatfactorn_hp'
+WVSAT = '0.0083556498*dvsatfactorn_hp'
+PVSAT = '-2.6650462e-11*dvsatfactorn_hp'
+A0 = 1.2529432
+LA0 = 2.2447635e-08
+WA0 = -3.4946308e-10
+PA0 = 8.4477928e-17
+AGS = -0.21154577
+LAGS = 1.245319e-07
+WAGS = 5.2192671e-08
+PAGS = -7.9748656e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.18606917
+LKETA = -1.867978e-08
+WKETA = -1.3940944e-08
+PKETA = 1.1962294e-15
+DWG = 0
+DWB = 0
+PCLM = 3.1003496
+LPCLM = -2.0493785e-07
+WPCLM = 3.1926064e-09
+PPCLM = -7.7145981e-16
+PDIBLC1 = 0
+PDIBLC2 = -0.060985236
+LPDIBLC2 = 1.1277245e-08
+WPDIBLC2 = 4.8019814e-09
+PPDIBLC2 = -7.3396758e-16
+PDIBLCB = -0.042878317
+LPDIBLCB = 2.1809914e-08
+WPDIBLCB = -3.3976507e-10
+PPDIBLCB = 8.2100616e-17
+DROUT = 0.56
+PVAG = 0.98362159
+LPVAG = -5.8558579e-08
+WPVAG = 9.1221398e-10
+PPVAG = -2.2043213e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.06158
+LPDITSD = -9.400132e-09
+WPDITSD = 1.4793296e-10
+PPDITSD = -3.5528101e-17
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -5.5747723e-11
+LALPHA0 = 3.9039053e-17
+WALPHA0 = -6.0814334e-19
+PALPHA0 = 1.4695475e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.026836199
+LAIGBINV = -5.8558416e-10
+WAIGBINV = 9.123929e-12
+PAIGBINV = -2.2044967e-18
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010144987
+LAIGC = 1.1613534e-11
+WAIGC = 1.3352312e-11
+PAIGC = -2.0672091e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5165257
+LUTE = 2.5781652e-08
+WUTE = 2.964158e-08
+PUTE = -4.5891341e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.610 NMOS
+LMIN = '1.33000000e-07+dlminn_hp'
+LMAX = '1.37000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.44427052+dvth0n610_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-7.3702402e-09+dlvth0n610_hp'
+WVTH0 = '-1.9970373e-08+dwvth0n610_hp'
+PVTH0 = '1.3170797e-15+dpvth0n610_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.16692634*dk2factorn_hp'
+LK2 = '8.6061702e-10*dk2factorn_hp'
+WK2 = '-1.3895874e-09*dk2factorn_hp'
+PK2 = '1.4631673e-17*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0.011853733
+LCDSCD = -1.721331e-09
+WCDSCD = 1.1910442e-10
+PCDSCD = -2.9256818e-17
+CIT = 0
+VOFF = -0.13330215
+LVOFF = -2.3018981e-09
+WVOFF = 3.9395551e-09
+PVOFF = -4.8516453e-17
+NFACTOR = 0.87389137
+LNFACTOR = 4.8210441e-08
+WNFACTOR = 3.8503461e-09
+PNFACTOR = -3.7973631e-16
+ETA0 = 0
+ETAB = -0.029807914
+LETAB = -6.298244e-09
+WETAB = 4.3579462e-10
+PETAB = -1.0704887e-16
+U0 = '(0.00481824*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.663611e-09*du0factorn_hp'
+WU0 = '1.9509607e-09*du0factorn_hp'
+PU0 = '-1.591153e-16*du0factorn_hp'
+UA = -3.1293525e-26
+LUA = 3.9224825e-33
+WUA = 2.7328529e-33
+PUA = -3.0149883e-40
+UB = 1e-19
+UC = -7.4912263e-28
+LUC = -5.0095984e-35
+WUC = 1.3706892e-34
+PUC = -1.4268602e-41
+EU = 2.9
+VSAT = '217091.59*dvsatfactorn_hp'
+LVSAT = '-0.021288442*dvsatfactorn_hp'
+WVSAT = '-0.0096896054*dvsatfactorn_hp'
+PVSAT = '2.3886908e-09*dvsatfactorn_hp'
+A0 = 1.2636812
+LA0 = 1.9795376e-08
+WA0 = -1.3695775e-09
+PA0 = 3.3644259e-16
+AGS = 1.1220182
+LAGS = -8.5373398e-08
+WAGS = -7.4495908e-08
+PAGS = 1.1966138e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.16747041
+LKETA = -1.7143987e-08
+WKETA = -1.2174063e-08
+PKETA = 1.0503291e-15
+DWG = 0
+DWB = 0
+PCLM = 3.002325
+LPCLM = -1.8072467e-07
+WPCLM = 1.2504945e-08
+PPCLM = -3.0717122e-15
+PDIBLC1 = 0
+PDIBLC2 = 0.061556861
+LPDIBLC2 = -8.0036491e-09
+WPDIBLC2 = -6.8395179e-09
+PPDIBLC2 = 1.0977174e-15
+PDIBLCB = -0.032446545
+LPDIBLCB = 1.9233119e-08
+WPDIBLCB = -1.3307834e-09
+PPDIBLCB = 3.2689621e-16
+DROUT = 0.56
+PVAG = 0.95561179
+LPVAG = -5.163991e-08
+WPVAG = 3.5731448e-09
+PPVAG = -8.777057e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.057101
+LPDITSD = -8.2912027e-09
+WPDITSD = 5.7334438e-10
+PPDITSD = -1.4087639e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -3.7074761e-11
+LALPHA0 = 3.4426627e-17
+WALPHA0 = -2.3820746e-18
+PALPHA0 = 5.8513522e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.026556159
+LAIGBINV = -5.1640293e-10
+WAIGBINV = 3.5727745e-11
+PAIGBINV = -8.7767134e-18
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010279297
+LAIGC = -8.6093995e-12
+WAIGC = 5.9285415e-13
+PAIGC = -1.460304e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5482057
+LUTE = 1.0844054e-08
+WUTE = 3.265118e-08
+PUTE = -3.1700623e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.011 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.32273358+dvth0n011_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0077024e-09+dlvth0n011_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14707612*dk2factorn_hp'
+LK2 = '1.1450578e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10204063
+LVOFF = -2.8060713e-10
+NFACTOR = 1.0594415
+LNFACTOR = 4.1773754e-08
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.035538061*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-5.7252892e-10*du0factorn_hp'
+UA = 3.4223936e-27
+LUA = -2.2855352e-34
+UB = 1e-19
+UC = -1.8852045e-27
+LUC = 1.5801795e-34
+EU = 2.9
+VSAT = '78678.208*dvsatfactorn_hp'
+LVSAT = '0.0018320923*dvsatfactorn_hp'
+A0 = 2.6863836
+LA0 = -1.1107059e-07
+AGS = 0.033910443
+LAGS = 9.1604612e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.1226133
+LPCLM = -5.9036193e-08
+PDIBLC1 = 0
+PDIBLC2 = -0.0051902983
+LPDIBLC2 = 2.8626441e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.45847762
+LPVAG = 2.2901152e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.3044778e-11
+LALPHA0 = 4.5802306e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027245673
+LAIGBINV = -6.870347e-10
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010347371
+LAIGC = -2.061113e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n011_hp'
+PVTH0 = '0.0+dpvth0n011_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.111 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.32429747+dvth0n111_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.1451548e-09+dlvth0n111_hp'
+WVTH0 = '-1.5526343e-08+dwvth0n111_hp'
+PVTH0 = '8.5633731e-15+dpvth0n111_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14646432*dk2factorn_hp'
+LK2 = '1.3846545e-09*dk2factorn_hp'
+WK2 = '-6.0739958e-09*dk2factorn_hp'
+PK2 = '-2.3787159e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.013883821
+LCDSCB = 1.4375799e-09
+WCDSCB = 8.8198572e-08
+PCDSCB = -1.4272293e-14
+CDSCD = -0.0059225471
+LCDSCD = 9.5838658e-10
+WCDSCD = 5.8799048e-08
+PCDSCD = -9.514862e-15
+CIT = 0
+VOFF = -0.098988039
+LVOFF = 5.5109077e-10
+WVOFF = -3.0306154e-08
+PVOFF = -8.2570967e-15
+NFACTOR = 1.115434
+LNFACTOR = 3.2685366e-08
+WNFACTOR = -5.5589297e-07
+PNFACTOR = 9.022952e-14
+ETA0 = 0
+ETAB = -0.073179195
+LETAB = -3.8381155e-14
+WETAB = -4.0186469e-12
+PETAB = 3.810481e-19
+U0 = '(0.035192265*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.5878378e-10*du0factorn_hp'
+WU0 = '3.4330577e-09*du0factorn_hp'
+PU0 = '8.5633834e-16*du0factorn_hp'
+UA = 3.4254055e-27
+LUA = -2.4867964e-34
+WUA = -2.99026e-35
+PUA = 1.9981218e-40
+UB = 1e-19
+UC = -1.9461279e-27
+LUC = 1.8760335e-34
+WUC = 6.0484759e-34
+PUC = -2.9372382e-40
+EU = 2.9
+VSAT = '79270.463*dvsatfactorn_hp'
+LVSAT = '0.0017362536*dvsatfactorn_hp'
+WVSAT = '-0.0058799065*dvsatfactorn_hp'
+PVSAT = '9.5148635e-10*dvsatfactorn_hp'
+A0 = 2.6863836
+LA0 = -1.1107059e-07
+AGS = 0.033910443
+LAGS = 9.1604612e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.1226133
+LPCLM = -5.9036193e-08
+PDIBLC1 = 0
+PDIBLC2 = -0.0051902983
+LPDIBLC2 = 2.8626441e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.34002669
+LPVAG = 4.2068882e-08
+WPVAG = 1.1759809e-06
+PPVAG = -1.9029723e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.3044778e-11
+LALPHA0 = 4.5802306e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027245673
+LAIGBINV = -6.870347e-10
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010335526
+LAIGC = -1.8694348e-11
+WAIGC = 1.17599e-10
+PAIGC = -1.9029809e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5226553
+LUTE = 5.8461533e-09
+WUTE = 6.1211358e-07
+PUTE = -5.804061e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.211 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.33842681+dvth0n211_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.6805153e-09+dlvth0n211_hp'
+WVTH0 = '-5.6911191e-08+dwvth0n211_hp'
+PVTH0 = '6.995302e-15+dpvth0n211_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14785792*dk2factorn_hp'
+LK2 = '8.3888804e-10*dk2factorn_hp'
+WK2 = '-1.9921355e-09*dk2factorn_hp'
+PK2 = '-7.8016588e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.022300431
+LCDSCB = -4.4253639e-09
+WCDSCB = -1.7785102e-08
+PCDSCB = 2.9002694e-15
+CDSCD = 0.014291114
+LCDSCD = -2.3254785e-09
+WCDSCD = -4.0676603e-10
+PCDSCD = 1.035789e-16
+CIT = 0
+VOFF = -0.12460531
+LVOFF = 2.8211786e-10
+WVOFF = 4.472682e-08
+PVOFF = -7.469275e-15
+NFACTOR = 1.1202659
+LNFACTOR = 4.1525346e-08
+WNFACTOR = -5.7004564e-07
+PNFACTOR = 6.4337216e-14
+ETA0 = 0
+ETAB = -0.096763452
+LETAB = 3.7691088e-09
+WETAB = 6.907427e-08
+PETAB = -1.1039451e-14
+U0 = '(0.042870128*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.1034284e-09*du0factorn_hp'
+WU0 = '-1.9055404e-08*du0factorn_hp'
+PU0 = '2.1587024e-15*du0factorn_hp'
+UA = 4.0702286e-27
+LUA = -2.6462347e-34
+WUA = -1.9185893e-33
+PUA = 2.4651165e-40
+UB = 1e-19
+UC = -3.5946097e-27
+LUC = 3.6262872e-34
+WUC = 5.4332509e-33
+PUC = -8.0637313e-40
+EU = 2.9
+VSAT = '75204.434*dvsatfactorn_hp'
+LVSAT = '0.0024019527*dvsatfactorn_hp'
+WVSAT = '0.0060294927*dvsatfactorn_hp'
+PVSAT = '-9.9834614e-10*dvsatfactorn_hp'
+A0 = 3.3589711
+LA0 = -1.7459009e-07
+WA0 = -1.9700086e-06
+PA0 = 1.860486e-13
+AGS = 0.028355416
+LAGS = 9.3019142e-08
+WAGS = 1.6270676e-08
+PAGS = -4.1431602e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.017109585
+LKETA = 2.0601462e-09
+WKETA = 3.7756026e-08
+PKETA = -6.0341682e-15
+DWG = 0
+DWB = 0
+PCLM = 2.1261933
+LPCLM = -5.994781e-08
+WPCLM = -1.0485889e-08
+PPCLM = 2.6701259e-15
+PDIBLC1 = 0
+PDIBLC2 = -0.008586497
+LPDIBLC2 = 3.4218847e-09
+WPDIBLC2 = 9.947466e-09
+PPDIBLC2 = -1.6380159e-15
+PDIBLCB = 0.035547923
+LPDIBLCB = 1.0300731e-08
+WPDIBLCB = 1.8878013e-07
+PPDIBLCB = -3.0170841e-14
+DROUT = 0.56
+PVAG = 0.61400697
+LPVAG = -2.6533211e-09
+WPVAG = 3.7349264e-07
+PPVAG = -5.9305896e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.96896
+LPDITSD = 4.9607876e-09
+WPDITSD = 9.0914993e-08
+PPDITSD = -1.4530147e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.5822288e-11
+LALPHA0 = 4.6509571e-17
+WALPHA0 = 8.1353268e-18
+PALPHA0 = -2.0715784e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027287336
+LAIGBINV = -6.9764368e-10
+WAIGBINV = -1.2203039e-10
+PAIGBINV = 3.107371e-17
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010383649
+LAIGC = -2.6610474e-11
+WAIGC = -2.3353699e-11
+PAIGC = 4.1565235e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.3128244
+LUTE = -1.4185402e-08
+WUTE = -2.4811588e-09
+PUTE = 6.3181582e-16
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.311 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29422383+dvth0n311_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.0546919e-08+dlvth0n311_hp'
+WVTH0 = '-1.5802416e-08+dwvth0n311_hp'
+PVTH0 = '6.0954654e-16+dpvth0n311_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.15624849*dk2factorn_hp'
+LK2 = '2.0511821e-09*dk2factorn_hp'
+WK2 = '5.811099e-09*dk2factorn_hp'
+PK2 = '-1.9075993e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0031002539
+LCDSCB = -1.2874132e-09
+WCDSCB = 7.1062828e-11
+PCDSCB = -1.8024819e-17
+CDSCD = 0.013724258
+LCDSCD = -2.1812638e-09
+WCDSCD = 1.2041002e-10
+PCDSCD = -3.0540795e-17
+CIT = 0
+VOFF = -0.067177449
+LVOFF = -8.5109414e-09
+WVOFF = -8.6810875e-09
+PVOFF = 7.0827011e-16
+NFACTOR = 0.27084404
+LNFACTOR = 1.481333e-07
+WNFACTOR = 2.1991668e-07
+PNFACTOR = -3.4808185e-14
+ETA0 = 0
+ETAB = -0.022963797
+LETAB = -7.9811077e-09
+WETAB = 4.4059069e-10
+PETAB = -1.1174977e-16
+U0 = '(0.018929107*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6685371e-09*du0factorn_hp'
+WU0 = '3.2097463e-09*du0factorn_hp'
+PU0 = '-4.1922556e-16*du0factorn_hp'
+UA = 2.0072553e-27
+LUA = 4.3623843e-37
+WUA = -2.4233504e-38
+PUA = 6.1226083e-45
+UB = 1e-19
+UC = 5.1749418e-28
+LUC = -2.2346628e-34
+WUC = 1.6089943e-33
+PUC = -2.6130478e-40
+EU = 2.9
+VSAT = '92697.899*dvsatfactorn_hp'
+LVSAT = '-0.00044939907*dvsatfactorn_hp'
+WVSAT = '-0.01023943*dvsatfactorn_hp'
+PVSAT = '1.653411e-09*dvsatfactorn_hp'
+A0 = 1.2421714
+LA0 = 2.5084492e-08
+WA0 = -1.3849082e-09
+PA0 = 3.5124227e-16
+AGS = 0.051029692
+LAGS = 8.7250549e-08
+WAGS = -4.8164016e-09
+PAGS = 1.2216319e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.0088598455
+LKETA = 3.4515025e-09
+WKETA = 4.5428284e-08
+PKETA = -7.3281295e-15
+DWG = 0
+DWB = 0
+PCLM = 1.1493723
+LPCLM = 9.8512178e-08
+WPCLM = 8.9795763e-07
+PPCLM = -1.4469766e-13
+PDIBLC1 = 0
+PDIBLC2 = 0.03669337
+LPDIBLC2 = -3.9101813e-09
+WPDIBLC2 = -3.2162811e-08
+PPDIBLC2 = 5.1808055e-15
+PDIBLCB = 0.4944393
+LPDIBLCB = -6.3175014e-08
+WPDIBLCB = -2.3798885e-07
+PPDIBLCB = 3.8161602e-14
+DROUT = 0.56
+PVAG = 1.0117278
+LPVAG = -6.5437915e-08
+WPVAG = 3.6123e-09
+PPVAG = -9.162234e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.066094
+LPDITSD = -1.0504766e-08
+WPDITSD = 5.8090104e-10
+PPDITSD = -1.4718192e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -7.4485151e-11
+LALPHA0 = 4.3625275e-17
+WALPHA0 = -2.4082113e-18
+PALPHA0 = 6.1081693e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027117279
+LAIGBINV = -6.5437929e-10
+WAIGBINV = 3.6122611e-11
+PAIGBINV = -9.1621742e-18
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010357241
+LAIGC = -2.1812565e-11
+WAIGC = 1.2053653e-12
+PAIGC = -3.0553211e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.2855579
+LUTE = -2.5222105e-08
+WUTE = -2.7839002e-08
+PUTE = 1.0895949e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.411 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26735463+dvth0n411_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.417776e-08+dlvth0n411_hp'
+WVTH0 = '-4.1949206e-09+dwvth0n411_hp'
+PVTH0 = '-9.5897667e-16+dpvth0n411_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13074114*dk2factorn_hp'
+LK2 = '-4.0216089e-09*dk2factorn_hp'
+WK2 = '-5.2080766e-09*dk2factorn_hp'
+PK2 = '7.1584639e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0090565847
+LCDSCB = -2.2605799e-09
+WCDSCB = -2.5020721e-09
+PCDSCB = 4.0238323e-16
+CDSCD = 0.014735151
+LCDSCD = -2.4332737e-09
+WCDSCD = -3.1629573e-10
+PCDSCD = 7.8327471e-17
+CIT = 0
+VOFF = -0.09330209
+LVOFF = -7.9315805e-09
+WVOFF = 2.6047578e-09
+PVOFF = 4.579862e-16
+NFACTOR = 0.93956446
+LNFACTOR = 4.5061569e-08
+WNFACTOR = -6.8970548e-08
+PNFACTOR = 9.7188049e-15
+ETA0 = 0
+ETAB = -0.019264946
+LETAB = -8.9032054e-09
+WETAB = -1.1573132e-09
+PETAB = 2.8659645e-16
+U0 = '(0.026181452*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '7.6828312e-10*du0factorn_hp'
+WU0 = '7.6733249e-11*du0factorn_hp'
+PU0 = '-3.0315828e-17*du0factorn_hp'
+UA = 2.9151476e-27
+LUA = -1.3919648e-34
+WUA = -3.9223371e-34
+PUA = 6.0327456e-41
+UB = 1e-19
+UC = 5.8308585e-27
+LUC = -1.1312772e-33
+WUC = -6.863791e-34
+PUC = 1.3086952e-40
+EU = 2.9
+VSAT = '65429.858*dvsatfactorn_hp'
+LVSAT = '0.0029514971*dvsatfactorn_hp'
+WVSAT = '0.0015403641*dvsatfactorn_hp'
+PVSAT = '1.8422382e-10*dvsatfactorn_hp'
+A0 = 1.2305456
+LA0 = 2.7982664e-08
+WA0 = 3.6374169e-09
+PA0 = -9.0076802e-16
+AGS = 0.010593987
+LAGS = 9.7330942e-08
+WAGS = 1.2651823e-08
+PAGS = -3.1330981e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.11841091
+LKETA = -1.4599642e-08
+WKETA = -1.8977741e-09
+PKETA = 4.6996479e-16
+DWG = 0
+DWB = 0
+PCLM = 3.3048489
+LPCLM = -2.5547245e-07
+WPCLM = -3.3208258e-08
+PPCLM = 8.2236969e-15
+PDIBLC1 = 0
+PDIBLC2 = -0.040385369
+LPDIBLC2 = 8.7331697e-09
+WPDIBLC2 = 1.1352046e-09
+PPDIBLC2 = -2.8112209e-16
+PDIBLCB = -0.064641584
+LPDIBLCB = 2.7187915e-08
+WPDIBLCB = 3.5340949e-09
+PPDIBLCB = -8.7518339e-16
+DROUT = 0.56
+PVAG = 1.0420546
+LPVAG = -7.2998211e-08
+WPVAG = -9.4888745e-09
+PPVAG = 2.3498243e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.070965
+LPDITSD = -1.1718766e-08
+WPDITSD = -1.5235353e-09
+PPDITSD = 3.7726583e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -9.4703043e-11
+LALPHA0 = 4.8665475e-17
+WALPHA0 = 6.325918e-18
+PALPHA0 = -1.5665498e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027420546
+LAIGBINV = -7.2998213e-10
+WAIGBINV = -9.4888855e-11
+PAIGBINV = 2.3498251e-17
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010458164
+LAIGC = -3.8301418e-11
+WAIGC = -4.2393215e-11
+PAIGC = 6.8176524e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.35
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.511 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.25492617+dvth0n511_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.1418773e-08+dlvth0n511_hp'
+WVTH0 = '-1.982655e-09+dwvth0n511_hp'
+PVTH0 = '-4.6787699e-16+dpvth0n511_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13533007*dk2factorn_hp'
+LK2 = '-1.1613449e-09*dk2factorn_hp'
+WK2 = '-4.3912475e-09*dk2factorn_hp'
+PK2 = '2.067194e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0.012787376
+LCDSCD = -1.9519517e-09
+WCDSCD = 3.04082e-11
+PCDSCD = -7.3478375e-18
+CIT = 0
+VOFF = -0.063600876
+LVOFF = -8.2727429e-09
+WVOFF = -2.6820584e-09
+PVOFF = 5.1871311e-16
+NFACTOR = 0.13737081
+LNFACTOR = 1.6312675e-07
+WNFACTOR = 7.3819923e-08
+PNFACTOR = -1.1296797e-14
+ETA0 = 0
+ETAB = -0.026391769
+LETAB = -7.1420723e-09
+WETAB = 1.112614e-10
+PETAB = -2.6885232e-17
+U0 = '(0.028052245*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-9.938434e-10*du0factorn_hp'
+WU0 = '-2.5626791e-10*du0factorn_hp'
+PU0 = '2.8334269e-16*du0factorn_hp'
+UA = 4.4180082e-27
+LUA = -4.2875346e-34
+WUA = -6.5974288e-34
+PUA = 1.118686e-40
+UB = 1e-19
+UC = 3.4411035e-27
+LUC = -6.2012179e-34
+WUC = -2.6100271e-34
+PUC = 3.9883863e-41
+EU = 2.9
+VSAT = '27141.884*dvsatfactorn_hp'
+LVSAT = '0.00413617*dvsatfactorn_hp'
+WVSAT = '0.0083556235*dvsatfactorn_hp'
+PVSAT = '-2.6647963e-11*dvsatfactorn_hp'
+A0 = 1.2529453
+LA0 = 2.2447439e-08
+WA0 = -3.4971584e-10
+PA0 = 8.4501896e-17
+AGS = -0.2115454
+LAGS = 1.2453186e-07
+WAGS = 5.2192635e-08
+PAGS = -7.9748621e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.18606916
+LKETA = -1.8679779e-08
+WKETA = -1.3940943e-08
+PKETA = 1.1962293e-15
+DWG = 0
+DWB = 0
+PCLM = 3.1003497
+LPCLM = -2.0493786e-07
+WPCLM = 3.1926063e-09
+PPCLM = -7.714598e-16
+PDIBLC1 = 0
+PDIBLC2 = -0.060985247
+LPDIBLC2 = 1.1277246e-08
+WPDIBLC2 = 4.8019829e-09
+PPDIBLC2 = -7.3396771e-16
+PDIBLCB = -0.042878333
+LPDIBLCB = 2.1809916e-08
+WPDIBLCB = -3.3976392e-10
+PPDIBLCB = 8.2100507e-17
+DROUT = 0.56
+PVAG = 0.98362129
+LPVAG = -5.8558551e-08
+WPVAG = 9.1224657e-10
+PPVAG = -2.2043522e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.061582
+LPDITSD = -9.4003823e-09
+WPDITSD = 1.4664931e-10
+PPDITSD = -3.5406385e-17
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -5.574753e-11
+LALPHA0 = 3.9039035e-17
+WALPHA0 = -6.0816329e-19
+PALPHA0 = 1.4695664e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.026836212
+LAIGBINV = -5.8558542e-10
+WAIGBINV = 9.1225108e-12
+PAIGBINV = -2.2043622e-18
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010144986
+LAIGC = 1.1613591e-11
+WAIGC = 1.3352418e-11
+PAIGC = -2.0672192e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5165279
+LUTE = 2.578186e-08
+WUTE = 2.9641971e-08
+PUTE = -4.5891711e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.611 NMOS
+LMIN = '1.37000000e-07+dlminn_hp'
+LMAX = '1.96000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.4442705+dvth0n611_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-7.3702381e-09+dlvth0n611_hp'
+WVTH0 = '-1.9970366e-08+dwvth0n611_hp'
+PVTH0 = '1.317079e-15+dpvth0n611_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.16692687*dk2factorn_hp'
+LK2 = '8.6066646e-10*dk2factorn_hp'
+WK2 = '-1.389552e-09*dk2factorn_hp'
+PK2 = '1.4628315e-17*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0.011853731
+LCDSCD = -1.7213308e-09
+WCDSCD = 1.1910448e-10
+PCDSCD = -2.9256824e-17
+CIT = 0
+VOFF = -0.13330216
+LVOFF = -2.3018969e-09
+WVOFF = 3.9395637e-09
+PVOFF = -4.8517268e-17
+NFACTOR = 0.87389878
+LNFACTOR = 4.8209739e-08
+WNFACTOR = 3.8497656e-09
+PNFACTOR = -3.7968126e-16
+ETA0 = 0
+ETAB = -0.029807938
+LETAB = -6.2982417e-09
+WETAB = 4.3579743e-10
+PETAB = -1.0704914e-16
+U0 = '(0.0048183235*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.6636031e-09*du0factorn_hp'
+WU0 = '1.9509546e-09*du0factorn_hp'
+PU0 = '-1.5911472e-16*du0factorn_hp'
+UA = -3.1293526e-26
+LUA = 3.9224827e-33
+WUA = 2.7328529e-33
+PUA = -3.0149883e-40
+UB = 1e-19
+UC = -7.4912944e-28
+LUC = -5.0095339e-35
+WUC = 1.3706942e-34
+PUC = -1.4268649e-41
+EU = 2.9
+VSAT = '217091.89*dvsatfactorn_hp'
+LVSAT = '-0.021288471*dvsatfactorn_hp'
+WVSAT = '-0.0096896272*dvsatfactorn_hp'
+PVSAT = '2.3886929e-09*dvsatfactorn_hp'
+A0 = 1.2636818
+LA0 = 1.9795327e-08
+WA0 = -1.3696827e-09
+PA0 = 3.3645257e-16
+AGS = 1.1220179
+LAGS = -8.5373369e-08
+WAGS = -7.449588e-08
+PAGS = 1.1966135e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.16747045
+LKETA = -1.7143991e-08
+WKETA = -1.2174066e-08
+PKETA = 1.0503294e-15
+DWG = 0
+DWB = 0
+PCLM = 3.0023256
+LPCLM = -1.8072473e-07
+WPCLM = 1.2504895e-08
+PPCLM = -3.0717075e-15
+PDIBLC1 = 0
+PDIBLC2 = 0.061556887
+LPDIBLC2 = -8.0036515e-09
+WPDIBLC2 = -6.8395198e-09
+PPDIBLC2 = 1.0977176e-15
+PDIBLCB = -0.032446342
+LPDIBLCB = 1.9233099e-08
+WPDIBLCB = -1.330803e-09
+PPDIBLCB = 3.2689807e-16
+DROUT = 0.56
+PVAG = 0.95561192
+LPVAG = -5.1639923e-08
+WPVAG = 3.5731358e-09
+PPVAG = -8.7770484e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.057093
+LPDITSD = -8.2904325e-09
+WPDITSD = 5.730832e-10
+PPDITSD = -1.4085162e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -3.7074557e-11
+LALPHA0 = 3.4426608e-17
+WALPHA0 = -2.3820957e-18
+PALPHA0 = 5.8513722e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.026556119
+LAIGBINV = -5.1639918e-10
+WAIGBINV = 3.5731348e-11
+PAIGBINV = -8.777055e-18
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010279267
+LAIGC = -8.6065114e-12
+WAIGC = 5.9579717e-13
+PAIGC = -1.4630946e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5481965
+LUTE = 1.0843181e-08
+WUTE = 3.2650487e-08
+PUTE = -3.1699966e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.012 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.32273357+dvth0n012_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0077038e-09+dlvth0n012_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14707595*dk2factorn_hp'
+LK2 = '1.1450322e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10204049
+LVOFF = -2.8062908e-10
+NFACTOR = 1.0594404
+LNFACTOR = 4.1773921e-08
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.035538056*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-5.7252824e-10*du0factorn_hp'
+UA = 3.4223908e-27
+LUA = -2.2855309e-34
+UB = 1e-19
+UC = -1.8852045e-27
+LUC = 1.5801797e-34
+EU = 2.9
+VSAT = '78678.237*dvsatfactorn_hp'
+LVSAT = '0.001832088*dvsatfactorn_hp'
+A0 = 2.6863837
+LA0 = -1.1107061e-07
+AGS = 0.033910652
+LAGS = 9.160458e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.1226153
+LPCLM = -5.9036494e-08
+PDIBLC1 = 0
+PDIBLC2 = -0.0051903191
+LPDIBLC2 = 2.8626473e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.45847737
+LPVAG = 2.290119e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.3044871e-11
+LALPHA0 = 4.580232e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027245652
+LAIGBINV = -6.8703146e-10
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010347365
+LAIGC = -2.0610216e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n012_hp'
+PVTH0 = '0.0+dpvth0n012_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.112 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.3242974+dvth0n112_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.1451649e-09+dlvth0n112_hp'
+WVTH0 = '-1.552578e-08+dwvth0n112_hp'
+PVTH0 = '8.5632864e-15+dpvth0n112_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14646403*dk2factorn_hp'
+LK2 = '1.3846108e-09*dk2factorn_hp'
+WK2 = '-6.0751614e-09*dk2factorn_hp'
+PK2 = '-2.3785366e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.013883821
+LCDSCB = 1.4375799e-09
+WCDSCB = 8.8198577e-08
+PCDSCB = -1.4272294e-14
+CDSCD = -0.0059225471
+LCDSCD = 9.5838658e-10
+WCDSCD = 5.8799048e-08
+PCDSCD = -9.5148619e-15
+CIT = 0
+VOFF = -0.098987783
+LVOFF = 5.5105136e-10
+WVOFF = -3.030728e-08
+PVOFF = -8.2569235e-15
+NFACTOR = 1.1154313
+LNFACTOR = 3.2685782e-08
+WNFACTOR = -5.558769e-07
+PNFACTOR = 9.0227048e-14
+ETA0 = 0
+ETAB = -0.073179197
+LETAB = -3.8096887e-14
+WETAB = -4.0002995e-12
+PETAB = 3.782259e-19
+U0 = '(0.035192254*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.5878214e-10*du0factorn_hp'
+WU0 = '3.4331207e-09*du0factorn_hp'
+PU0 = '8.5632864e-16*du0factorn_hp'
+UA = 3.4254008e-27
+LUA = -2.4867891e-34
+WUA = -2.9883102e-35
+PUA = 1.9980918e-40
+UB = 1e-19
+UC = -1.9461279e-27
+LUC = 1.8760335e-34
+WUC = 6.0484664e-34
+PUC = -2.9372367e-40
+EU = 2.9
+VSAT = '79270.494*dvsatfactorn_hp'
+LVSAT = '0.0017362489*dvsatfactorn_hp'
+WVSAT = '-0.005879932*dvsatfactorn_hp'
+PVSAT = '9.5149028e-10*dvsatfactorn_hp'
+A0 = 2.6863837
+LA0 = -1.1107061e-07
+AGS = 0.033910652
+LAGS = 9.160458e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.1226153
+LPCLM = -5.9036494e-08
+PDIBLC1 = 0
+PDIBLC2 = -0.0051903191
+LPDIBLC2 = 2.8626473e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.34002623
+LPVAG = 4.2068953e-08
+WPVAG = 1.175983e-06
+PPVAG = -1.9029755e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.3044871e-11
+LALPHA0 = 4.580232e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027245652
+LAIGBINV = -6.8703146e-10
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010335532
+LAIGC = -1.8695212e-11
+WAIGC = 1.1748422e-10
+PAIGC = -1.9012155e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5226565
+LUTE = 5.8463483e-09
+WUTE = 6.1212617e-07
+PUTE = -5.8042546e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.212 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.33842699+dvth0n212_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.6804874e-09+dlvth0n212_hp'
+WVTH0 = '-5.6911352e-08+dwvth0n212_hp'
+PVTH0 = '6.9953267e-15+dpvth0n212_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14785809*dk2factorn_hp'
+LK2 = '8.3891373e-10*dk2factorn_hp'
+WK2 = '-1.9919801e-09*dk2factorn_hp'
+PK2 = '-7.8018977e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.022300434
+LCDSCB = -4.4253643e-09
+WCDSCB = -1.7785106e-08
+PCDSCB = 2.9002699e-15
+CDSCD = 0.014291114
+LCDSCD = -2.3254785e-09
+WCDSCD = -4.0676611e-10
+PCDSCD = 1.0357892e-16
+CIT = 0
+VOFF = -0.12460563
+LVOFF = 2.8216725e-10
+WVOFF = 4.4727385e-08
+PVOFF = -7.4693619e-15
+NFACTOR = 1.1202703
+LNFACTOR = 4.1524668e-08
+WNFACTOR = -5.7005043e-07
+PNFACTOR = 6.4337952e-14
+ETA0 = 0
+ETAB = -0.096763435
+LETAB = 3.7691062e-09
+WETAB = 6.9074233e-08
+PETAB = -1.1039445e-14
+U0 = '(0.042870143*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.1034307e-09*du0factorn_hp'
+WU0 = '-1.9055416e-08*du0factorn_hp'
+PU0 = '2.1587042e-15*du0factorn_hp'
+UA = 4.070232e-27
+LUA = -2.64624e-34
+WUA = -1.9185938e-33
+PUA = 2.4651235e-40
+UB = 1e-19
+UC = -3.5946109e-27
+LUC = 3.626289e-34
+WUC = 5.4332534e-33
+PUC = -8.0637352e-40
+EU = 2.9
+VSAT = '75204.462*dvsatfactorn_hp'
+LVSAT = '0.0024019484*dvsatfactorn_hp'
+WVSAT = '0.0060294758*dvsatfactorn_hp'
+PVSAT = '-9.9834354e-10*dvsatfactorn_hp'
+A0 = 3.3589718
+LA0 = -1.745902e-07
+WA0 = -1.9700104e-06
+PA0 = 1.8604888e-13
+AGS = 0.028355772
+LAGS = 9.3019088e-08
+WAGS = 1.6270244e-08
+PAGS = -4.1430938e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.017109573
+LKETA = 2.0601479e-09
+WKETA = 3.7756059e-08
+PKETA = -6.0341733e-15
+DWG = 0
+DWB = 0
+PCLM = 2.1261958
+LPCLM = -5.9948196e-08
+WPCLM = -1.0487515e-08
+PPCLM = 2.6703761e-15
+PDIBLC1 = 0
+PDIBLC2 = -0.0085865228
+LPDIBLC2 = 3.4218887e-09
+WPDIBLC2 = 9.9474805e-09
+PPDIBLC2 = -1.6380181e-15
+PDIBLCB = 0.035547922
+LPDIBLCB = 1.0300731e-08
+WPDIBLCB = 1.8878014e-07
+PPDIBLCB = -3.0170842e-14
+DROUT = 0.56
+PVAG = 0.61400735
+LPVAG = -2.6533805e-09
+WPVAG = 3.7349224e-07
+PPVAG = -5.9305835e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.96896
+LPDITSD = 4.9608577e-09
+WPDITSD = 9.0916328e-08
+PPDITSD = -1.4530352e-14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.5822311e-11
+LALPHA0 = 4.6509574e-17
+WALPHA0 = 8.135122e-18
+PALPHA0 = -2.0715469e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027287307
+LAIGBINV = -6.9763929e-10
+WAIGBINV = -1.2200829e-10
+PAIGBINV = 3.1070309e-17
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010383604
+LAIGC = -2.6603606e-11
+WAIGC = -2.332123e-11
+PAIGC = 4.1515292e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.3128213
+LUTE = -1.4185872e-08
+WUTE = -2.4812273e-09
+PUTE = 6.3182636e-16
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.312 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29422398+dvth0n312_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.0546896e-08+dlvth0n312_hp'
+WVTH0 = '-1.580255e-08+dwvth0n312_hp'
+PVTH0 = '6.0956716e-16+dpvth0n312_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.15624869*dk2factorn_hp'
+LK2 = '2.0512118e-09*dk2factorn_hp'
+WK2 = '5.8112786e-09*dk2factorn_hp'
+PK2 = '-1.907627e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0031002508
+LCDSCB = -1.2874127e-09
+WCDSCB = 7.1064473e-11
+PCDSCB = -1.8025072e-17
+CDSCD = 0.013724258
+LCDSCD = -2.1812638e-09
+WCDSCD = 1.2040995e-10
+PCDSCD = -3.0540783e-17
+CIT = 0
+VOFF = -0.0671768
+LVOFF = -8.5110412e-09
+WVOFF = -8.6814244e-09
+PVOFF = 7.0832193e-16
+NFACTOR = 0.27084119
+LNFACTOR = 1.4813374e-07
+WNFACTOR = 2.1991865e-07
+PNFACTOR = -3.4808488e-14
+ETA0 = 0
+ETAB = -0.022963815
+LETAB = -7.9811049e-09
+WETAB = 4.4058625e-10
+PETAB = -1.1174908e-16
+U0 = '(0.018929109*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6685368e-09*du0factorn_hp'
+WU0 = '3.2097461e-09*du0factorn_hp'
+PU0 = '-4.1922553e-16*du0factorn_hp'
+UA = 2.0072522e-27
+LUA = 4.3671709e-37
+WUA = -2.2626026e-38
+PUA = 5.8753461e-45
+UB = 1e-19
+UC = 5.1749805e-28
+LUC = -2.2346687e-34
+WUC = 1.6089921e-33
+PUC = -2.6130445e-40
+EU = 2.9
+VSAT = '92697.906*dvsatfactorn_hp'
+LVSAT = '-0.00044940007*dvsatfactorn_hp'
+WVSAT = '-0.010239427*dvsatfactorn_hp'
+PVSAT = '1.6534105e-09*dvsatfactorn_hp'
+A0 = 1.2421689
+LA0 = 2.508488e-08
+WA0 = -1.3836707e-09
+PA0 = 3.5105193e-16
+AGS = 0.05102958
+LAGS = 8.7250566e-08
+WAGS = -4.8163982e-09
+PAGS = 1.2216313e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.0088598788
+LKETA = 3.4514973e-09
+WKETA = 4.5428275e-08
+PKETA = -7.3281282e-15
+DWG = 0
+DWB = 0
+PCLM = 1.149374
+LPCLM = 9.8511922e-08
+WPCLM = 8.9795679e-07
+PPCLM = -1.4469753e-13
+PDIBLC1 = 0
+PDIBLC2 = 0.036693369
+LPDIBLC2 = -3.910181e-09
+WPDIBLC2 = -3.2162819e-08
+PPDIBLC2 = 5.1808067e-15
+PDIBLCB = 0.49443951
+LPDIBLCB = -6.3175046e-08
+WPDIBLCB = -2.3798904e-07
+PPDIBLCB = 3.8161631e-14
+DROUT = 0.56
+PVAG = 1.0117278
+LPVAG = -6.5437922e-08
+WPVAG = 3.6122211e-09
+PPVAG = -9.1621126e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.066097
+LPDITSD = -1.0505238e-08
+WPDITSD = 5.7896198e-10
+PPDITSD = -1.4688365e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -7.4485574e-11
+LALPHA0 = 4.362534e-17
+WALPHA0 = -2.408044e-18
+PALPHA0 = 6.1079119e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027117285
+LAIGBINV = -6.543802e-10
+WAIGBINV = 3.6112661e-11
+PAIGBINV = -9.1606438e-18
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010357246
+LAIGC = -2.1813188e-11
+WAIGC = 1.1925415e-12
+PAIGC = -3.0355955e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.2855523
+LUTE = -2.522296e-08
+WUTE = -2.7841405e-08
+PUTE = 1.0896319e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.412 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.24737608+dvth0n412_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.7250859e-08+dlvth0n412_hp'
+WVTH0 = '4.435742e-09+dwvth0n412_hp'
+PVTH0 = '-2.2865452e-15+dpvth0n412_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1169746*dk2factorn_hp'
+LK2 = '-6.1391789e-09*dk2factorn_hp'
+WK2 = '-1.1155128e-08*dk2factorn_hp'
+PK2 = '1.6306218e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0090565859
+LCDSCB = -2.2605801e-09
+WCDSCB = -2.5020723e-09
+PCDSCB = 4.0238326e-16
+CDSCD = 0.0238161
+LCDSCD = -3.8301053e-09
+WCDSCD = -4.2392659e-09
+PCDSCD = 6.8175874e-16
+CIT = 0
+VOFF = -0.068888997
+LVOFF = -1.1686803e-08
+WVOFF = -7.9417553e-09
+PVOFF = 2.0802509e-15
+NFACTOR = 0.48551984
+LNFACTOR = 1.1490271e-07
+WNFACTOR = 1.2717747e-07
+PNFACTOR = -2.0452683e-14
+ETA0 = 0
+ETAB = 0.013961646
+LETAB = -1.401412e-08
+WETAB = -1.5511213e-08
+PETAB = 2.4945133e-15
+U0 = '(0.021621709*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.4696628e-09*du0factorn_hp'
+WU0 = '2.046543e-09*du0factorn_hp'
+PU0 = '-3.3331196e-16*du0factorn_hp'
+UA = 2.0052375e-27
+LUA = 7.6589422e-37
+WUA = 8.4772118e-37
+PUA = -1.3632917e-43
+UB = 1e-19
+UC = 7.6352412e-27
+LUC = -1.4088273e-33
+WUC = -1.4658729e-33
+PUC = 2.5077126e-40
+EU = 2.9
+VSAT = '47267.986*dvsatfactorn_hp'
+LVSAT = '0.0057451563*dvsatfactorn_hp'
+WVSAT = '0.0093862985*dvsatfactorn_hp'
+PVSAT = '-1.0226378e-09*dvsatfactorn_hp'
+A0 = 1.1261153
+LA0 = 4.4046143e-08
+WA0 = 4.8751482e-08
+PA0 = -7.8402134e-15
+AGS = -0.35264417
+LAGS = 1.5320424e-07
+WAGS = 1.6957066e-07
+PAGS = -2.7270354e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.17289663
+LKETA = -2.2980635e-08
+WKETA = -2.54356e-08
+PKETA = 4.0905531e-15
+DWG = 0
+DWB = 0
+PCLM = 4.2156608
+LPCLM = -3.9557353e-07
+WPCLM = -4.2667911e-07
+PPCLM = 6.8747383e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.068388799
+LPDIBLC2 = 1.3040657e-08
+WPDIBLC2 = 1.3232678e-08
+PPDIBLC2 = -2.1419554e-15
+PDIBLCB = -0.16610696
+LPDIBLCB = 4.279532e-08
+WPDIBLCB = 4.736704e-08
+PPDIBLCB = -7.617567e-15
+DROUT = 0.56
+PVAG = 1.2285828
+LPVAG = -1.0168998e-07
+WPVAG = -9.0069133e-08
+PPVAG = 1.474468e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.114696
+LPDITSD = -1.8445458e-08
+WPDITSD = -2.0415914e-08
+PPDITSD = 3.2832915e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -4.5986932e-10
+LALPHA0 = 1.0483535e-16
+WALPHA0 = 1.6407773e-16
+PALPHA0 = -2.5831934e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.030144802
+LAIGBINV = -1.1490271e-09
+WAIGBINV = -1.2717747e-09
+PAIGBINV = 2.0452683e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010494839
+LAIGC = -4.394277e-11
+WAIGC = -5.82479e-11
+PAIGC = 9.25642e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.35
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.512 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30505363+dvth0n512_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.7081666e-09+dlvth0n512_hp'
+WVTH0 = '-5.8308614e-09+dwvth0n512_hp'
+PVTH0 = '1.2405412e-16+dpvth0n512_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.18876424*dk2factorn_hp'
+LK2 = '7.0578984e-09*dk2factorn_hp'
+WK2 = '1.6234277e-09*dk2factorn_hp'
+PK2 = '-7.1845794e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = -0.0037506294
+LCDSCD = 5.9192433e-10
+WCDSCD = 6.6761203e-10
+PCDSCD = -1.0536253e-16
+CIT = 0
+VOFF = -0.127261
+LVOFF = 1.5194576e-09
+WVOFF = 2.4484614e-09
+PVOFF = -2.7046345e-16
+NFACTOR = 1.2817178
+LNFACTOR = -1.2896703e-08
+WNFACTOR = -1.4545769e-08
+PNFACTOR = 2.2956132e-15
+ETA0 = 0
+ETAB = -0.086903318
+LETAB = 2.165814e-09
+WETAB = 2.4427506e-09
+PETAB = -3.8551489e-16
+U0 = '(0.035978377*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.2130411e-09*du0factorn_hp'
+WU0 = '-5.0894403e-10*du0factorn_hp'
+PU0 = '3.2220933e-16*du0factorn_hp'
+UA = 3.7550179e-27
+LUA = -3.2677229e-34
+WUA = -3.1061318e-34
+PUA = 5.8165468e-41
+UB = 1e-19
+UC = -1.4246453e-27
+LUC = 1.2832769e-34
+WUC = 1.4678686e-34
+PUC = -2.2842328e-41
+EU = 2.9
+VSAT = '61342.857*dvsatfactorn_hp'
+LVSAT = '-0.0011246237*dvsatfactorn_hp'
+WVSAT = '0.0068809715*dvsatfactorn_hp'
+PVSAT = '2.0018301e-10*dvsatfactorn_hp'
+A0 = 1.4431301
+LA0 = -6.8067864e-09
+WA0 = -7.6771511e-09
+PA0 = 1.211608e-15
+AGS = 0.67501259
+LAGS = -1.1838487e-08
+WAGS = -1.3352242e-08
+PAGS = 2.1072508e-15
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.030362538
+LKETA = 5.2710131e-09
+WKETA = -6.4531714e-11
+PKETA = -9.3824033e-16
+DWG = 0
+DWB = 0
+PCLM = 1.4416491
+LPCLM = 5.0203455e-08
+WPCLM = 6.7094966e-08
+PPCLM = -1.0600921e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.010701831
+LPDIBLC2 = 2.5033996e-10
+WPDIBLC2 = -8.4545425e-10
+PPDIBLC2 = 1.3472106e-16
+PDIBLCB = 0.14190733
+LPDIBLCB = -6.6138152e-09
+WPDIBLCB = -7.4595052e-09
+PPDIBLCB = 1.1772591e-15
+DROUT = 0.56
+PVAG = 0.64401239
+LPVAG = -6.3199104e-09
+WPVAG = 1.3984398e-08
+PPVAG = -2.2311936e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.981954
+LPDITSD = 2.8480278e-09
+WPDITSD = 3.2121971e-09
+PPDITSD = -5.0694895e-16
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 6.0948219e-10
+LALPHA0 = -6.3286601e-17
+WALPHA0 = -2.6266835e-17
+PALPHA0 = 4.0937735e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.021874807
+LAIGBINV = 1.7757801e-10
+WAIGBINV = 2.0028441e-10
+PAIGBINV = -3.1608885e-17
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010134312
+LAIGC = 1.3255504e-11
+WAIGC = 5.9259037e-12
+PAIGC = -9.2487272e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.3916336
+LUTE = 6.5706085e-09
+WUTE = 7.4107738e-09
+PUTE = -1.1695683e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.612 NMOS
+LMIN = '1.96000000e-07+dlminn_hp'
+LMAX = '2.00000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.48082635+dvth0n612_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.299326e-08+dlvth0n612_hp'
+WVTH0 = '-2.252927e-08+dwvth0n612_hp'
+PVTH0 = '1.7106897e-15+dpvth0n612_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12938945*dk2factorn_hp'
+LK2 = '-4.9133395e-09*dk2factorn_hp'
+WK2 = '-4.0171774e-09*dk2factorn_hp'
+PK2 = '4.1880966e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = -0.025502538
+LCDSCD = 4.0248105e-09
+WCDSCD = 2.7340433e-09
+PCDSCD = -4.3148672e-16
+CIT = 0
+VOFF = -0.16998982
+LVOFF = 3.341399e-09
+WVOFF = 6.5076993e-09
+PVOFF = -4.4354789e-16
+NFACTOR = 1.6877878
+LNFACTOR = -7.6982676e-08
+WNFACTOR = -5.3122421e-08
+PNFACTOR = 8.3837806e-15
+ETA0 = 0
+ETAB = -0.1664922
+LETAB = 1.4726532e-08
+WETAB = 1.0003695e-08
+PETAB = -1.5787831e-15
+U0 = '(0.024830555*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '5.8532163e-10*du0factorn_hp'
+WU0 = '5.5009909e-10*du0factorn_hp'
+PU0 = '5.6364874e-17*du0factorn_hp'
+UA = -1.9847697e-26
+LUA = 2.1618853e-33
+WUA = 1.9316448e-33
+PUA = -1.78257e-40
+UB = 1e-19
+UC = -2.9273913e-27
+LUC = 2.849649e-34
+WUC = 2.8954773e-34
+PUC = -3.7722864e-41
+EU = 2.9
+VSAT = '288068.99*dvsatfactorn_hp'
+LVSAT = '-0.032206169*dvsatfactorn_hp'
+WVSAT = '-0.014658012*dvsatfactorn_hp'
+PVSAT = '3.1529298e-09*dvsatfactorn_hp'
+A0 = 1.6932863
+LA0 = -4.6286442e-08
+WA0 = -3.1441992e-08
+PA0 = 4.9621752e-15
+AGS = 1.8691433
+LAGS = -2.0029619e-07
+WAGS = -1.2679466e-07
+PAGS = 2.0010733e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.13084172
+LKETA = -1.150976e-08
+WKETA = -9.6100541e-09
+PKETA = 6.559331e-16
+DWG = 0
+DWB = 0
+PCLM = -0.74464528
+LPCLM = 3.9563433e-07
+WPCLM = 2.7479294e-07
+PPCLM = -4.3416854e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.10807029
+LPDIBLC2 = -1.5158343e-08
+WPDIBLC2 = -1.0095458e-08
+PPDIBLC2 = 1.5985459e-15
+PDIBLCB = 0.38494924
+LPDIBLCB = -4.4970689e-08
+WPDIBLCB = -3.0548487e-08
+PPDIBLCB = 4.8211622e-15
+DROUT = 0.56
+PVAG = 0.18798447
+LPVAG = 6.6436533e-08
+WPVAG = 5.7307051e-08
+PPVAG = -9.1430557e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.877082
+LPDITSD = 1.939885e-08
+WPDITSD = 1.3174991e-08
+PPDITSD = -2.079277e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.4644509e-09
+LALPHA0 = -1.9653805e-16
+WALPHA0 = -1.0748887e-16
+PALPHA0 = 1.6752661e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.015349224
+LAIGBINV = 1.2074455e-09
+WAIGBINV = 8.2021477e-10
+PAIGBINV = -1.294463e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0099417008
+LAIGC = 4.3317867e-11
+WAIGC = 2.4223984e-11
+PAIGC = -3.7807972e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.9628481
+LUTE = 7.4624881e-08
+WUTE = 6.1676152e-08
+PUTE = -7.6347242e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.013 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.3227337+dvth0n013_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0076824e-09+dlvth0n013_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14707625*dk2factorn_hp'
+LK2 = '1.1450795e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10204065
+LVOFF = -2.8060353e-10
+NFACTOR = 1.0594409
+LNFACTOR = 4.1773852e-08
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.035538048*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-5.7252696e-10*du0factorn_hp'
+UA = 3.4223943e-27
+LUA = -2.2855365e-34
+UB = 1e-19
+UC = -1.8852045e-27
+LUC = 1.5801797e-34
+EU = 2.9
+VSAT = '78678.19*dvsatfactorn_hp'
+LVSAT = '0.0018320952*dvsatfactorn_hp'
+A0 = 2.6863829
+LA0 = -1.1107047e-07
+AGS = 0.033910313
+LAGS = 9.1604633e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.1226116
+LPCLM = -5.9035917e-08
+PDIBLC1 = 0
+PDIBLC2 = -0.0051902805
+LPDIBLC2 = 2.8626412e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.45847768
+LPVAG = 2.2901142e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.3044646e-11
+LALPHA0 = 4.5802285e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027245674
+LAIGBINV = -6.8703491e-10
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010347361
+LAIGC = -2.0609515e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n013_hp'
+PVTH0 = '0.0+dpvth0n013_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.113 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.3242977+dvth0n113_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.145118e-09+dlvth0n113_hp'
+WVTH0 = '-1.552738e-08+dwvth0n113_hp'
+PVTH0 = '8.5635389e-15+dpvth0n113_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14646456*dk2factorn_hp'
+LK2 = '1.384694e-09*dk2factorn_hp'
+WK2 = '-6.0729002e-09*dk2factorn_hp'
+PK2 = '-2.3788935e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.01388382
+LCDSCB = 1.4375797e-09
+WCDSCB = 8.8198564e-08
+PCDSCB = -1.4272292e-14
+CDSCD = -0.0059225471
+LCDSCD = 9.5838657e-10
+WCDSCD = 5.8799047e-08
+PCDSCD = -9.5148618e-15
+CIT = 0
+VOFF = -0.098988095
+LVOFF = 5.5110057e-10
+WVOFF = -3.0305793e-08
+PVOFF = -8.2571583e-15
+NFACTOR = 1.1154334
+LNFACTOR = 3.2685438e-08
+WNFACTOR = -5.5589416e-07
+PNFACTOR = 9.0229773e-14
+ETA0 = 0
+ETAB = -0.073179201
+LETAB = -3.7406378e-14
+WETAB = -3.9568615e-12
+PETAB = 3.7137052e-19
+U0 = '(0.035192246*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.5878073e-10*du0factorn_hp'
+WU0 = '3.4331288e-09*du0factorn_hp'
+PU0 = '8.5632737e-16*du0factorn_hp'
+UA = 3.4254069e-27
+LUA = -2.4867988e-34
+WUA = -2.9908953e-35
+PUA = 1.9981326e-40
+UB = 1e-19
+UC = -1.9461275e-27
+LUC = 1.8760328e-34
+WUC = 6.0484265e-34
+PUC = -2.9372305e-40
+EU = 2.9
+VSAT = '79270.44*dvsatfactorn_hp'
+LVSAT = '0.0017362574*dvsatfactorn_hp'
+WVSAT = '-0.0058798529*dvsatfactorn_hp'
+PVSAT = '9.514778e-10*dvsatfactorn_hp'
+A0 = 2.6863829
+LA0 = -1.1107047e-07
+AGS = 0.033910313
+LAGS = 9.1604633e-08
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.1226116
+LPCLM = -5.9035917e-08
+PDIBLC1 = 0
+PDIBLC2 = -0.0051902805
+LPDIBLC2 = 2.8626412e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.34002679
+LPVAG = 4.2068865e-08
+WPVAG = 1.1759804e-06
+PPVAG = -1.9029715e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -8.3044646e-11
+LALPHA0 = 4.5802285e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.027245674
+LAIGBINV = -6.8703491e-10
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010335506
+LAIGC = -1.8691102e-11
+WAIGC = 1.1769869e-10
+PAIGC = -1.9046002e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5226549
+LUTE = 5.8460825e-09
+WUTE = 6.1210945e-07
+PUTE = -5.8039907e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.213 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.32380092+dvth0n213_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '5.988775e-09+dlvth0n213_hp'
+WVTH0 = '-1.4072299e-08+dwvth0n213_hp'
+PVTH0 = '2.3446744e-16+dpvth0n213_hp'
+K1 = '0.64076895*dk1factorn_hp'
+LK1 = '1.7724838e-09*dk1factorn_hp'
+WK1 = '3.2895736e-08*dk1factorn_hp'
+PK1 = '-5.191605e-15*dk1factorn_hp'
+K2 = '-0.14005831*dk2factorn_hp'
+LK2 = '-3.9204678e-10*dk2factorn_hp'
+WK2 = '-2.4836804e-08*dk2factorn_hp'
+PK2 = '2.8251804e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.024202453
+LCDSCB = -4.725541e-09
+WCDSCB = -2.335613e-08
+PCDSCB = 3.779489e-15
+CDSCD = 0.017513718
+LCDSCD = -2.8340698e-09
+WCDSCD = -9.8457723e-09
+PCDSCD = 1.5932429e-15
+CIT = 0
+VOFF = -0.10708651
+LVOFF = -2.4826996e-09
+WVOFF = -6.5855312e-09
+PVOFF = 6.2884254e-16
+NFACTOR = 1.02153
+LNFACTOR = 5.7107862e-08
+WNFACTOR = -2.8085098e-07
+PNFACTOR = 1.8696495e-14
+ETA0 = 0
+ETAB = -0.084972367
+LETAB = 1.9082399e-09
+WETAB = 3.4538226e-08
+PETAB = -5.5889729e-15
+U0 = '(0.040473749*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.2523169e-10*du0factorn_hp'
+WU0 = '-1.2036394e-08*du0factorn_hp'
+PU0 = '1.0509622e-15*du0factorn_hp'
+UA = 3.7014517e-27
+LUA = -2.064231e-34
+WUA = -8.3844427e-34
+PUA = 7.6043141e-41
+UB = 1e-19
+UC = -2.1794887e-27
+LUC = 1.3929432e-34
+WUC = 1.2883578e-33
+PUC = -1.5222609e-40
+EU = 2.9
+VSAT = '70151.112*dvsatfactorn_hp'
+LVSAT = '0.0031994681*dvsatfactorn_hp'
+WVSAT = '0.020830658*dvsatfactorn_hp'
+PVSAT = '-3.3342662e-09*dvsatfactorn_hp'
+A0 = 3.0723309
+LA0 = -1.2935254e-07
+WA0 = -1.1304419e-06
+PA0 = 5.3548187e-14
+AGS = -0.10054888
+LAGS = 1.1336282e-07
+WAGS = 3.9383098e-07
+PAGS = -6.3729729e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.0235548
+LKETA = 1.0429623e-09
+WKETA = 1.8877992e-08
+PKETA = -3.0548367e-15
+DWG = 0
+DWB = 0
+PCLM = 2.1946246
+LPCLM = -7.0747623e-08
+WPCLM = -2.1092606e-07
+PPCLM = 3.4303587e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.0094435357
+LPDIBLC2 = 3.5571425e-09
+WPDIBLC2 = 1.2457784e-08
+PPDIBLC2 = -2.0341943e-15
+PDIBLCB = 0.067773961
+LPDIBLCB = 5.2148176e-09
+WPDIBLCB = 9.4390068e-08
+PPDIBLCB = -1.5274201e-14
+DROUT = 0.56
+PVAG = 0.68146733
+LPVAG = -1.3299914e-08
+WPVAG = 1.7590108e-07
+PPVAG = -2.8121999e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 13.984471
+LPDITSD = 2.5128974e-09
+WPDITSD = 4.5484344e-08
+PPDITSD = -7.3602766e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -2.126692e-10
+LALPHA0 = 6.652855e-17
+WALPHA0 = 3.7967031e-16
+PALPHA0 = -6.0707231e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.02825412
+LAIGBINV = -8.5022175e-10
+WAIGBINV = -2.9537404e-09
+PAIGBINV = 4.7797427e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010428367
+LAIGC = -3.3668009e-11
+WAIGC = -1.5429214e-10
+PAIGC = 2.4821358e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.2551056
+LUTE = -2.329457e-08
+WUTE = -1.7154242e-07
+PUTE = 2.7313064e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.313 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.34556661+dvth0n313_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.4440026e-09+dlvth0n313_hp'
+WVTH0 = '-3.431439e-08+dwvth0n313_hp'
+PVTH0 = '3.5311058e-15+dpvth0n313_hp'
+K1 = '0.69708205*dk1factorn_hp'
+LK1 = '-7.1148496e-09*dk1factorn_hp'
+WK1 = '-1.9475447e-08*dk1factorn_hp'
+PK1 = '3.073615e-15*dk1factorn_hp'
+K2 = '-0.18582699*dk2factorn_hp'
+LK2 = '6.71926e-09*dk2factorn_hp'
+WK2 = '1.772807e-08*dk2factorn_hp'
+PK2 = '-3.7883349e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.0027422234
+LCDSCB = -3.6535341e-10
+WCDSCB = 1.7024193e-09
+PCDSCB = -2.7548549e-16
+CDSCD = 0.0038253374
+LCDSCD = -6.1901609e-10
+WCDSCD = 2.8844214e-09
+PCDSCD = -4.6675708e-16
+CIT = 0
+VOFF = -0.13407234
+LVOFF = 2.0464123e-09
+WVOFF = 1.8511285e-08
+PVOFF = -3.5832315e-15
+NFACTOR = 0.5071572
+LNFACTOR = 1.1083835e-07
+WNFACTOR = 1.9751573e-07
+PNFACTOR = -3.127286e-14
+ETA0 = 0
+ETAB = -0.059182602
+LETAB = -2.265056e-09
+WETAB = 1.0553744e-08
+PETAB = -1.7078077e-15
+U0 = '(0.027548548*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.0821688e-10*du0factorn_hp'
+WU0 = '-1.5957839e-11*du0factorn_hp'
+PU0 = '8.9855067e-17*du0factorn_hp'
+UA = 2.3831934e-27
+LUA = -5.8894325e-35
+WUA = 3.8753595e-34
+PUA = -6.1158619e-41
+UB = 1e-19
+UC = -3.6421538e-27
+LUC = 4.3300938e-34
+WUC = 2.6486363e-33
+PUC = -4.253811e-40
+EU = 2.9
+VSAT = '96747.211*dvsatfactorn_hp'
+LVSAT = '-0.0010884615*dvsatfactorn_hp'
+WVSAT = '-0.0039037136*dvsatfactorn_hp'
+PVSAT = '6.5350825e-10*dvsatfactorn_hp'
+A0 = 2.1242369
+LA0 = -1.1412309e-07
+WA0 = -2.4871446e-07
+PA0 = 3.9384797e-14
+AGS = 0.44698641
+LAGS = 2.4760659e-08
+WAGS = -1.1537684e-07
+PAGS = 1.8670281e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.0012091508
+LKETA = 4.6589352e-09
+WKETA = 3.9659445e-08
+PKETA = -6.4176915e-15
+DWG = 0
+DWB = 0
+PCLM = 1.1798065
+LPCLM = 9.370907e-08
+WPCLM = 7.328548e-07
+PPCLM = -1.1864114e-13
+PDIBLC1 = 0
+PDIBLC2 = 0.030694394
+LPDIBLC2 = -2.9634228e-09
+WPDIBLC2 = -2.487049e-08
+PPDIBLC2 = 4.0299315e-15
+PDIBLCB = 0.3311508
+LPDIBLCB = -3.7404823e-08
+WPDIBLCB = -1.505504e-07
+PPDIBLCB = 2.4362065e-14
+DROUT = 0.56
+PVAG = 0.80469497
+LPVAG = -3.2764e-08
+WPVAG = 6.1299376e-08
+PPVAG = -1.0020398e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.018456
+LPDITSD = -2.986612e-09
+WPDITSD = 1.3877968e-08
+PPDITSD = -2.2457328e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.1555118e-10
+LALPHA0 = -1.793026e-17
+WALPHA0 = -1.1157464e-16
+PALPHA0 = 1.7839463e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.024147587
+LAIGBINV = -1.8570248e-10
+WAIGBINV = 8.6533588e-10
+PAIGBINV = -1.4002865e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010219872
+LAIGC = -1.32846e-13
+WAIGC = 3.9608357e-11
+PAIGC = -6.3663435e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5172502
+LUTE = 1.1343602e-08
+WUTE = 7.2252088e-08
+PUTE = -4.9004363e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.413 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26181754+dvth0n413_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.4971709e-08+dlvth0n413_hp'
+WVTH0 = '1.8652081e-09+dwvth0n413_hp'
+PVTH0 = '-1.8808635e-15+dpvth0n413_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12036468*dk2factorn_hp'
+LK2 = '-5.6041566e-09*dk2factorn_hp'
+WK2 = '-1.0551651e-08*dk2factorn_hp'
+PK2 = '1.5353811e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = 0.0055424361
+LCDSCB = -1.705977e-09
+WCDSCB = -1.8765536e-09
+PCDSCB = 3.0366391e-16
+CDSCD = 0.017862075
+LCDSCD = -2.8904411e-09
+WCDSCD = -3.1794494e-09
+PCDSCD = 5.1449851e-16
+CIT = 0
+VOFF = -0.075606168
+LVOFF = -1.0626699e-08
+WVOFF = -6.7460988e-09
+PVOFF = 1.8915523e-15
+NFACTOR = 0.79924267
+LNFACTOR = 6.5390975e-08
+WNFACTOR = 7.1334804e-08
+PNFACTOR = -1.1639594e-14
+ETA0 = 0
+ETAB = -0.0078232267
+LETAB = -1.0576031e-08
+WETAB = -1.1633506e-08
+PETAB = 1.8825335e-15
+U0 = '(0.023581898*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.1603058e-09*du0factorn_hp'
+WU0 = '1.6976353e-09*du0factorn_hp'
+PU0 = '-2.7824735e-16*du0factorn_hp'
+UA = 4.1704548e-27
+LUA = -3.4094869e-34
+WUA = -3.8456095e-34
+PUA = 6.0688867e-41
+UB = 1e-19
+UC = 4.6536452e-27
+LUC = -9.3827183e-34
+WUC = -9.3514884e-34
+PUC = 1.6701239e-40
+EU = 2.9
+VSAT = '79098.746*dvsatfactorn_hp'
+LVSAT = '0.00072162561*dvsatfactorn_hp'
+WVSAT = '0.0037204231*dvsatfactorn_hp'
+PVSAT = '-1.2844936e-10*dvsatfactorn_hp'
+A0 = 1.6525822
+LA0 = -3.9040863e-08
+WA0 = -4.4959626e-08
+PA0 = 6.9492736e-15
+AGS = -0.11448313
+LAGS = 1.1561766e-07
+WAGS = 1.27178e-07
+PAGS = -2.0579943e-14
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.13717244
+LKETA = -1.7342644e-08
+WKETA = -1.9076694e-08
+PKETA = 3.0869905e-15
+DWG = 0
+DWB = 0
+PCLM = 3.6174154
+LPCLM = -3.0115845e-07
+WPCLM = -3.2019227e-07
+PPCLM = 5.1941631e-14
+PDIBLC1 = 0
+PDIBLC2 = -0.049881836
+LPDIBLC2 = 1.0119888e-08
+WPDIBLC2 = 9.9384412e-09
+PPDIBLC2 = -1.622059e-15
+PDIBLCB = -0.099579719
+LPDIBLCB = 3.229599e-08
+WPDIBLCB = 3.552519e-08
+PPDIBLCB = -5.7486862e-15
+DROUT = 0.56
+PVAG = 1.1035785
+LPVAG = -8.19618e-08
+WPVAG = -6.7818289e-08
+PPVAG = 1.1233052e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14.086028
+LPDITSD = -1.392106e-08
+WPDITSD = -1.5312994e-08
+PPDITSD = 2.4779486e-15
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = -2.2628957e-10
+LALPHA0 = 6.7971797e-17
+WALPHA0 = 1.2250057e-16
+PALPHA0 = -1.9270226e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.028358635
+LAIGBINV = -8.6713435e-10
+WAIGBINV = -9.5383706e-10
+PAIGBINV = 1.5434991e-16
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010412429
+LAIGC = -3.0936795e-11
+WAIGC = -4.357639e-11
+PAIGC = 6.9409622e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.35
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.513 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30138384+dvth0n513_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.2873336e-09+dlvth0n513_hp'
+WVTH0 = '-5.1775935e-09+dwvth0n513_hp'
+PVTH0 = '2.0955368e-17+dpvth0n513_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.19253296*dk2factorn_hp'
+LK2 = '7.6526782e-09*dk2factorn_hp'
+WK2 = '2.2943034e-09*dk2factorn_hp'
+PK2 = '-8.2433554e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.12357771
+LVOFF = 9.3816047e-10
+WVOFF = 1.7928355e-09
+PVOFF = -1.6699256e-16
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.07318
+U0 = '(0.033969143*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.8959437e-09*du0factorn_hp'
+WU0 = '-1.5129435e-10*du0factorn_hp'
+PU0 = '2.6576506e-16*du0factorn_hp'
+UA = 2.6058446e-27
+LUA = -1.4540976e-34
+WUA = -1.0606033e-34
+PUA = 2.5882937e-41
+UB = 1e-19
+UC = -1.2059449e-27
+LUC = 9.3812393e-35
+WUC = 1.0785819e-34
+PUC = -1.6698606e-41
+EU = 2.9
+VSAT = '54216.867*dvsatfactorn_hp'
+WVSAT = '0.0081493976*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.034040118
+LKETA = 4.6906174e-09
+WKETA = -7.1914098e-10
+PKETA = -8.3492989e-16
+DWG = 0
+DWB = 0
+PCLM = 1.8178379
+LPCLM = -9.1666511e-09
+WPCLM = 1.3253192e-10
+PPCLM = -3.2909424e-17
+PDIBLC1 = 0
+PDIBLC2 = 0.0060318449
+LPDIBLC2 = 9.873571e-10
+WPDIBLC2 = -1.4194076e-11
+PPDIBLC2 = 3.5315844e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72108472
+LPVAG = -1.8483466e-08
+WPVAG = 2.6559468e-10
+PPVAG = -6.6092009e-17
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.5872662e-10
+LALPHA0 = -3.9494357e-17
+WALPHA0 = 5.6768468e-19
+PALPHA0 = -1.4125037e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010168268
+LAIGC = 7.8966064e-12
+WAIGC = -1.1572348e-13
+PAIGC = 2.861689e-20
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.35
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.613 NMOS
+LMIN = '2.00000000e-07+dlminn_hp'
+LMAX = '2.04000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.43525933+dvth0n613_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.8018721e-09+dlvth0n613_hp'
+WVTH0 = '-1.7895765e-08+dwvth0n613_hp'
+PVTH0 = '9.7942991e-16+dpvth0n613_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13585311*dk2factorn_hp'
+LK2 = '-3.8932446e-09*dk2factorn_hp'
+WK2 = '-3.0902826e-09*dk2factorn_hp'
+PK2 = '2.7252712e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 1.9164184e-16
+LCDSCD = -3.1011483e-23
+WCDSCD = -1.8205975e-23
+PCDSCD = 2.9460909e-30
+CIT = 0
+VOFF = -0.21104876
+LVOFF = 9.8213201e-09
+WVOFF = 1.0102585e-08
+PVOFF = -1.0108927e-15
+NFACTOR = 2.690312
+LNFACTOR = -2.3520105e-07
+WNFACTOR = -1.4157964e-07
+PNFACTOR = 2.2344099e-14
+ETA0 = 0
+ETAB = -0.07318
+U0 = '(-0.015523656*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '6.9540232e-09*du0factorn_hp'
+WU0 = '4.5505215e-09*du0factorn_hp'
+PU0 = '-5.7498179e-16*du0factorn_hp'
+UA = -9.1336923e-27
+LUA = 4.7100097e-34
+WUA = 1.0091957e-33
+PUA = -3.2676082e-41
+UB = 1e-19
+UC = 8.5173711e-28
+LUC = -3.1145714e-34
+WUC = -8.7621598e-35
+PUC = 2.1802e-41
+EU = 2.9
+VSAT = '121258.08*dvsatfactorn_hp'
+LVSAT = '-0.0058800708*dvsatfactorn_hp'
+WVSAT = '0.001780482*dvsatfactorn_hp'
+PVSAT = '5.5860673e-10*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.066959317
+LKETA = 1.97072e-08
+WKETA = 8.8758053e-09
+PKETA = -2.2615052e-15
+DWG = 0
+DWB = 0
+PCLM = 1.8183122
+LPCLM = -8.8516207e-09
+WPCLM = 8.747011e-11
+PPCLM = -6.2837313e-17
+PDIBLC1 = 0
+PDIBLC2 = 0.0059820632
+LPDIBLC2 = 9.5322071e-10
+WPDIBLC2 = -9.4648107e-12
+PPDIBLC2 = 6.7745417e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.7220136
+LPVAG = -1.7843945e-08
+WPVAG = 1.7735123e-10
+PPVAG = -1.2684646e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.607148e-10
+LALPHA0 = -3.8128407e-17
+WALPHA0 = 3.7880765e-19
+PALPHA0 = -2.7101563e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010167858
+LAIGC = 7.6257759e-12
+WAIGC = -7.675696e-14
+PAIGC = 5.4345784e-20
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.49
+WUTE = 1.33e-08
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.014 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.32499766+dvth0n014_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.6413282e-09+dlvth0n014_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11406887
+LVOFF = 1.6658025e-09
+NFACTOR = 1.3186967
+LNFACTOR = -1.7892049e-10
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.032*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 4.1726948e-27
+LUA = -3.4996728e-34
+UB = 1e-19
+UC = -6.6539685e-28
+LUC = -3.9371315e-35
+EU = 2.9
+VSAT = '90000*dvsatfactorn_hp'
+A0 = 1.7296631
+LA0 = 4.3745921e-08
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8212189
+LPCLM = -1.0264557e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0057415798
+LPDIBLC2 = 1.0936476e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72659089
+LPVAG = -2.0484938e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7033684e-10
+LALPHA0 = -4.3745907e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165932
+LAIGC = 8.7493323e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n014_hp'
+PVTH0 = '0.0+dpvth0n014_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.114 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.31634829+dvth0n114_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.4314923e-09+dlvth0n114_hp'
+WVTH0 = '8.5871013e-08+dwvth0n114_hp'
+PVTH0 = '-7.8447491e-15+dpvth0n114_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13507924*dk2factorn_hp'
+LK2 = '-4.57678e-10*dk2factorn_hp'
+WK2 = '-4.8853277e-08*dk2factorn_hp'
+PK2 = '4.5438271e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10831849
+LVOFF = 2.0609456e-09
+WVOFF = -5.7089738e-08
+PVOFF = -3.9229802e-15
+NFACTOR = 1.3189882
+LNFACTOR = -2.5379663e-10
+WNFACTOR = -2.8945163e-09
+PNFACTOR = 7.4337034e-16
+ETA0 = 0
+ETAB = -0.073179885
+LETAB = 7.3210506e-14
+WETAB = 2.8297188e-12
+PETAB = -7.268339e-19
+U0 = '(0.032365635*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0137867e-10*du0factorn_hp'
+WU0 = '-3.630028e-09*du0factorn_hp'
+PU0 = '1.9992874e-15*du0factorn_hp'
+UA = 3.7119348e-27
+LUA = -2.9504582e-34
+WUA = 4.574426e-33
+PUA = -5.4526022e-40
+UB = 1e-19
+UC = 2.3712523e-28
+LUC = -1.6569066e-34
+WUC = -8.9602392e-33
+PUC = 1.2540985e-39
+EU = 2.9
+VSAT = '84343.358*dvsatfactorn_hp'
+LVSAT = '0.00091535773*dvsatfactorn_hp'
+WVSAT = '0.056159137*dvsatfactorn_hp'
+PVSAT = '-9.0876716e-09*dvsatfactorn_hp'
+A0 = 1.8427958
+LA0 = 2.5438782e-08
+WA0 = -1.1231818e-06
+PA0 = 1.8175328e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8212189
+LPCLM = -1.0264557e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0057415798
+LPDIBLC2 = 1.0936476e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72659089
+LPVAG = -2.0484938e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7033684e-10
+LALPHA0 = -4.3745907e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165932
+LAIGC = 8.7493323e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4175167
+LUTE = -1.1167372e-08
+WUTE = -4.3170203e-07
+PUTE = 1.1086967e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.214 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.34825202+dvth0n214_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0320982e-09+dlvth0n214_hp'
+WVTH0 = '-7.5750101e-09+dwvth0n214_hp'
+PVTH0 = '-8.1692388e-16+dpvth0n214_hp'
+K1 = '0.62953779*dk1factorn_hp'
+LK1 = '3.5899111e-09*dk1factorn_hp'
+WK1 = '6.5791822e-08*dk1factorn_hp'
+PK1 = '-1.051485e-14*dk1factorn_hp'
+K2 = '-0.13697772*dk2factorn_hp'
+LK2 = '-8.9054763e-10*dk2factorn_hp'
+WK2 = '-4.3292631e-08*dk2factorn_hp'
+PK2 = '5.8117023e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11663785
+LVOFF = -9.371015e-10
+WVOFF = -3.2722332e-08
+PVOFF = 4.8582997e-15
+NFACTOR = 1.4976875
+LNFACTOR = -1.9943948e-08
+WNFACTOR = -5.2630475e-07
+PNFACTOR = 5.8415825e-14
+ETA0 = 0
+ETAB = -0.073178916
+LETAB = -1.7644755e-13
+WETAB = -9.5659177e-15
+PETAB = 4.4145435e-21
+U0 = '(0.030402383*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '9.0451667e-10*du0factorn_hp'
+WU0 = '2.120337e-09*du0factorn_hp'
+PU0 = '-1.23988e-15*du0factorn_hp'
+UA = 6.0558261e-27
+LUA = -5.8740795e-34
+WUA = -2.2908317e-33
+PUA = 3.1106847e-40
+UB = 1e-19
+UC = -2.3503261e-27
+LUC = 1.6693923e-34
+WUC = -1.3815942e-33
+PUC = 2.7982554e-40
+EU = 2.9
+VSAT = '103565.82*dvsatfactorn_hp'
+LVSAT = '-0.0022076992*dvsatfactorn_hp'
+WVSAT = '-0.00014343859*dvsatfactorn_hp'
+PVSAT = '5.9762197e-11*dvsatfactorn_hp'
+A0 = 0.98776665
+LA0 = 2.0797165e-07
+WA0 = 1.3811986e-06
+PA0 = -3.5288549e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8214489
+LPCLM = -1.0360327e-08
+WPCLM = -6.7346786e-10
+PPCLM = 2.805127e-16
+PDIBLC1 = 0
+PDIBLC2 = 0.0057170934
+LPDIBLC2 = 1.1038495e-09
+WPDIBLC2 = 7.1720563e-11
+PPDIBLC2 = -2.9881414e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72704953
+LPVAG = -2.0676026e-08
+WPVAG = -1.3433456e-09
+PPVAG = 5.5969474e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7131628e-10
+LALPHA0 = -4.415398e-17
+WALPHA0 = -2.8687718e-18
+PALPHA0 = 1.1952439e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165736
+LAIGC = 8.8309356e-12
+WAIGC = 5.7360077e-13
+PAIGC = -2.39016e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5655032
+LUTE = 2.6933968e-08
+WUTE = 1.7502522e-09
+PUTE = -7.2915645e-16
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.314 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.38217867+dvth0n314_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-3.4805621e-09+dlvth0n314_hp'
+WVTH0 = '-3.9126802e-08+dwvth0n314_hp'
+PVTH0 = '4.3098502e-15+dpvth0n314_hp'
+K1 = '0.74216459*dk1factorn_hp'
+LK1 = '-1.4410105e-08*dk1factorn_hp'
+WK1 = '-3.8951101e-08*dk1factorn_hp'
+PK1 = '6.2251654e-15*dk1factorn_hp'
+K2 = '-0.21194816*dk2factorn_hp'
+LK2 = '1.0946188e-08*dk2factorn_hp'
+WK2 = '2.6429879e-08*dk2factorn_hp'
+PK2 = '-5.1964617e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.19411369
+LVOFF = 1.1762304e-08
+WVOFF = 3.9330196e-08
+PVOFF = -6.9521477e-15
+NFACTOR = 0.42344242
+LNFACTOR = 1.2438508e-07
+WNFACTOR = 4.7274319e-07
+PNFACTOR = -7.5810167e-14
+ETA0 = 0
+ETAB = -0.073178928
+LETAB = -1.7049632e-13
+WETAB = 2.0814072e-15
+PETAB = -1.1201001e-21
+U0 = '(0.034168318*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.6299419e-10*du0factorn_hp'
+WU0 = '-1.3819818e-09*du0factorn_hp'
+PU0 = '3.1090507e-16*du0factorn_hp'
+UA = 5.5043145e-28
+LUA = 2.3768322e-34
+WUA = 2.8291853e-33
+PUA = -4.5626632e-40
+UB = 1e-19
+UC = -4.7603301e-27
+LUC = 6.1395268e-34
+WUC = 8.597095e-34
+PUC = -1.3589696e-40
+EU = 2.9
+VSAT = '68326.54*dvsatfactorn_hp'
+LVSAT = '0.0035105716*dvsatfactorn_hp'
+WVSAT = '0.032629088*dvsatfactorn_hp'
+PVSAT = '-5.2582297e-09*dvsatfactorn_hp'
+A0 = 2.469274
+LA0 = -1.6995699e-07
+WA0 = 3.3968114e-09
+PA0 = -1.4118488e-15
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8205105
+LPCLM = -9.9696548e-09
+WPCLM = 1.9922456e-10
+PPCLM = -8.2812734e-17
+PDIBLC1 = 0
+PDIBLC2 = 0.0058170424
+LPDIBLC2 = 1.0622302e-09
+WPDIBLC2 = -2.1232048e-11
+PPDIBLC2 = 8.824522e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72517748
+LPVAG = -1.9896481e-08
+WPVAG = 3.9765753e-10
+PPVAG = -1.6528197e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.6731846e-10
+LALPHA0 = -4.2489242e-17
+WALPHA0 = 8.4919882e-19
+PALPHA0 = -3.5296221e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010166535
+LAIGC = 8.4980514e-12
+WAIGC = -1.6985251e-13
+PAIGC = 7.0566307e-20
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7489311
+LUTE = 4.8834204e-08
+WUTE = 1.7233823e-07
+PUTE = -2.1096376e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.414 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30514045+dvth0n414_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '7.9611956e-09+dlvth0n414_hp'
+WVTH0 = '-5.8462889e-09+dwvth0n414_hp'
+PVTH0 = '-6.3298909e-16+dpvth0n414_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1305321*dk2factorn_hp'
+LK2 = '-3.9588648e-09*dk2factorn_hp'
+WK2 = '-8.7418618e-09*dk2factorn_hp'
+PK2 = '1.242521e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.095759532
+LVOFF = -7.3654814e-09
+WVOFF = -3.1588002e-09
+PVOFF = 1.3110557e-15
+NFACTOR = 1.7404343
+LNFACTOR = -8.6912656e-08
+WNFACTOR = -9.6197308e-08
+PNFACTOR = 1.5470453e-14
+ETA0 = 0
+ETAB = -0.073178169
+LETAB = -2.9438784e-13
+WETAB = -3.2594216e-13
+PETAB = 5.2401035e-20
+U0 = '(0.029462682*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.0867723e-10*du0factorn_hp'
+WU0 = '6.5085267e-10*du0factorn_hp'
+PU0 = '-1.0885699e-16*du0factorn_hp'
+UA = 1.0666109e-26
+LUA = -1.3920755e-33
+WUA = -1.5407874e-33
+PUA = 2.4778943e-40
+UB = 1e-19
+UC = -4.291154e-27
+LUC = 5.0917556e-34
+WUC = 6.5702541e-34
+PUC = -9.063325e-41
+EU = 2.9
+VSAT = '174591.15*dvsatfactorn_hp'
+LVSAT = '-0.014730956*dvsatfactorn_hp'
+WVSAT = '-0.013277225*dvsatfactorn_hp'
+PVSAT = '2.6221101e-09*dvsatfactorn_hp'
+A0 = 3.231981
+LA0 = -2.9461918e-07
+WA0 = -3.2609261e-07
+PA0 = 5.2442213e-14
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8226438
+LPCLM = -1.0728503e-08
+WPCLM = -7.2236284e-10
+PPCLM = 2.4500987e-16
+PDIBLC1 = 0
+PDIBLC2 = 0.0056388007
+LPDIBLC2 = 1.135539e-09
+WPDIBLC2 = 5.576837e-11
+PPDIBLC2 = -2.284489e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72856574
+LPVAG = -2.1277243e-08
+WPVAG = -1.0660693e-09
+PPVAG = 4.3120728e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7444788e-10
+LALPHA0 = -4.5421538e-17
+WALPHA0 = -2.2307123e-18
+PALPHA0 = 9.1378998e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165108
+LAIGC = 9.0846474e-12
+WAIGC = 4.4663255e-13
+PAIGC = -1.8284318e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.35
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.514 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30138372+dvth0n514_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.2873528e-09+dlvth0n514_hp'
+WVTH0 = '-5.1775907e-09+dwvth0n514_hp'
+PVTH0 = '2.0954918e-17+dpvth0n514_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.19253305*dk2factorn_hp'
+LK2 = '7.6526924e-09*dk2factorn_hp'
+WK2 = '2.2943072e-09*dk2factorn_hp'
+PK2 = '-8.2433617e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.12357748
+LVOFF = 9.3812315e-10
+WVOFF = 1.7927944e-09
+PVOFF = -1.6698592e-16
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.07318
+U0 = '(0.033969128*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.8959413e-09*du0factorn_hp'
+WU0 = '-1.5129465e-10*du0factorn_hp'
+PU0 = '2.6576511e-16*du0factorn_hp'
+UA = 2.6058406e-27
+LUA = -1.4540911e-34
+WUA = -1.0605962e-34
+PUA = 2.5882822e-41
+UB = 1e-19
+UC = -1.2059446e-27
+LUC = 9.3812346e-35
+WUC = 1.0785814e-34
+PUC = -1.6698598e-41
+EU = 2.9
+VSAT = '54216.867*dvsatfactorn_hp'
+WVSAT = '0.0081493976*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.034040118
+LKETA = 4.6906174e-09
+WKETA = -7.1914099e-10
+PKETA = -8.3492989e-16
+DWG = 0
+DWB = 0
+PCLM = 1.8178454
+LPCLM = -9.167861e-09
+WPCLM = 1.3175987e-10
+PPCLM = -3.278449e-17
+PDIBLC1 = 0
+PDIBLC2 = 0.0060318362
+LPDIBLC2 = 9.8735852e-10
+WPDIBLC2 = -1.4191944e-11
+PPDIBLC2 = 3.5312394e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72108405
+LPVAG = -1.8483356e-08
+WPVAG = 2.6567215e-10
+PPVAG = -6.6104545e-17
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.5872661e-10
+LALPHA0 = -3.9494355e-17
+WALPHA0 = 5.6767396e-19
+PALPHA0 = -1.4124863e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010168256
+LAIGC = 7.8985235e-12
+WAIGC = -1.136841e-13
+PAIGC = 2.8286877e-20
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.35
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.614 NMOS
+LMIN = '2.04000000e-07+dlminn_hp'
+LMAX = '2.91000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.43525951+dvth0n614_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.8019009e-09+dlvth0n614_hp'
+WVTH0 = '-1.7895791e-08+dwvth0n614_hp'
+PVTH0 = '9.7943402e-16+dpvth0n614_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13585329*dk2factorn_hp'
+LK2 = '-3.8932155e-09*dk2factorn_hp'
+WK2 = '-3.09027e-09*dk2factorn_hp'
+PK2 = '2.7252508e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.21104955
+LVOFF = 9.8214483e-09
+WVOFF = 1.0102641e-08
+PVOFF = -1.0109018e-15
+NFACTOR = 2.6903068
+LNFACTOR = -2.3520019e-07
+WNFACTOR = -1.4157914e-07
+PNFACTOR = 2.2344018e-14
+ETA0 = 0
+ETAB = -0.07318
+U0 = '(-0.015523708*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '6.9540317e-09*du0factorn_hp'
+WU0 = '4.5505248e-09*du0factorn_hp'
+PU0 = '-5.7498232e-16*du0factorn_hp'
+UA = -9.1336755e-27
+LUA = 4.7099825e-34
+WUA = 1.0091944e-33
+PUA = -3.2675877e-41
+UB = 1e-19
+UC = 8.5173616e-28
+LUC = -3.1145699e-34
+WUC = -8.7621531e-35
+PUC = 2.1801989e-41
+EU = 2.9
+VSAT = '121257.68*dvsatfactorn_hp'
+LVSAT = '-0.0058800049*dvsatfactorn_hp'
+WVSAT = '0.0017805207*dvsatfactorn_hp'
+PVSAT = '5.5860046e-10*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.066959296
+LKETA = 1.9707196e-08
+WKETA = 8.8758033e-09
+PKETA = -2.2615049e-15
+DWG = 0
+DWB = 0
+PCLM = 1.8183062
+LPCLM = -8.8506496e-09
+WPCLM = 8.7978436e-11
+PPCLM = -6.291957e-17
+PDIBLC1 = 0
+PDIBLC2 = 0.0059821404
+LPDIBLC2 = 9.5320821e-10
+WPDIBLC2 = -9.4708449e-12
+PPDIBLC2 = 6.7755181e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72201432
+LPVAG = -1.7844062e-08
+WPVAG = 1.7729608e-10
+PPVAG = -1.2683753e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.6071443e-10
+LALPHA0 = -3.8128346e-17
+WALPHA0 = 3.7883151e-19
+PALPHA0 = -2.7101949e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010167856
+LAIGC = 7.6261041e-12
+WAIGC = -7.56504e-14
+PAIGC = 5.4166721e-20
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.49
+WUTE = 1.33e-08
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.015 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.3249982+dvth0n015_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.6411955e-09+dlvth0n015_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11406873
+LVOFF = 1.6657687e-09
+NFACTOR = 1.3186981
+LNFACTOR = -1.7928402e-10
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.032*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 4.1726942e-27
+LUA = -3.4996712e-34
+UB = 1e-19
+UC = -6.6539652e-28
+LUC = -3.9371399e-35
+EU = 2.9
+VSAT = '90000*dvsatfactorn_hp'
+A0 = 1.7296656
+LA0 = 4.37453e-08
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8212136
+LPCLM = -1.0263224e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0057415771
+LPDIBLC2 = 1.0936482e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72659085
+LPVAG = -2.0484929e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7033693e-10
+LALPHA0 = -4.3745929e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165953
+LAIGC = 8.7440275e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n015_hp'
+PVTH0 = '0.0+dpvth0n015_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.115 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.31634908+dvth0n115_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.4312958e-09+dlvth0n115_hp'
+WVTH0 = '8.5868471e-08+dwvth0n115_hp'
+PVTH0 = '-7.8441165e-15+dpvth0n115_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135079*dk2factorn_hp'
+LK2 = '-4.5773828e-10*dk2factorn_hp'
+WK2 = '-4.8855682e-08*dk2factorn_hp'
+PK2 = '4.5444256e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10831812
+LVOFF = 2.0608518e-09
+WVOFF = -5.7092131e-08
+PVOFF = -3.9223849e-15
+NFACTOR = 1.3189903
+LNFACTOR = -2.5431229e-10
+WNFACTOR = -2.9005864e-09
+PNFACTOR = 7.448807e-16
+ETA0 = 0
+ETAB = -0.073179882
+LETAB = 7.2395702e-14
+WETAB = 2.7972078e-12
+PETAB = -7.1874453e-19
+U0 = '(0.032365635*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0137852e-10*du0factorn_hp'
+WU0 = '-3.6300221e-09*du0factorn_hp'
+PU0 = '1.9992859e-15*du0factorn_hp'
+UA = 3.7119345e-27
+LUA = -2.9504576e-34
+WUA = 4.5744219e-33
+PUA = -5.452592e-40
+UB = 1e-19
+UC = 2.3712753e-28
+LUC = -1.6569124e-34
+WUC = -8.9602587e-33
+PUC = 1.2541034e-39
+EU = 2.9
+VSAT = '84343.357*dvsatfactorn_hp'
+LVSAT = '0.0009153581*dvsatfactorn_hp'
+WVSAT = '0.056159152*dvsatfactorn_hp'
+PVSAT = '-9.0876752e-09*dvsatfactorn_hp'
+A0 = 1.8428
+LA0 = 2.5437743e-08
+WA0 = -1.1231985e-06
+PA0 = 1.8175742e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8212136
+LPCLM = -1.0263224e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0057415771
+LPDIBLC2 = 1.0936482e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72659085
+LPVAG = -2.0484929e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7033693e-10
+LALPHA0 = -4.3745929e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165953
+LAIGC = 8.7440275e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4175167
+LUTE = -1.1167366e-08
+WUTE = -4.3170181e-07
+PUTE = 1.1086961e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.215 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.34825165+dvth0n215_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0321894e-09+dlvth0n215_hp'
+WVTH0 = '-7.5741674e-09+dwvth0n215_hp'
+PVTH0 = '-8.1713357e-16+dpvth0n215_hp'
+K1 = '0.62953766*dk1factorn_hp'
+LK1 = '3.5899428e-09*dk1factorn_hp'
+WK1 = '6.5792195e-08*dk1factorn_hp'
+PK1 = '-1.0514942e-14*dk1factorn_hp'
+K2 = '-0.13697866*dk2factorn_hp'
+LK2 = '-8.9031469e-10*dk2factorn_hp'
+WK2 = '-4.3291585e-08*dk2factorn_hp'
+PK2 = '5.8114419e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11663839
+LVOFF = -9.3696711e-10
+WVOFF = -3.2722038e-08
+PVOFF = 4.8582266e-15
+NFACTOR = 1.4976886
+LNFACTOR = -1.9944208e-08
+WNFACTOR = -5.2630781e-07
+PNFACTOR = 5.8416585e-14
+ETA0 = 0
+ETAB = -0.07317893
+LETAB = -1.7299335e-13
+WETAB = 8.1759992e-15
+PETAB = -2.9740378e-28
+U0 = '(0.030402375*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '9.0451874e-10*du0factorn_hp'
+WU0 = '2.1203656e-09*du0factorn_hp'
+PU0 = '-1.2398871e-15*du0factorn_hp'
+UA = 6.0558237e-27
+LUA = -5.8740737e-34
+WUA = -2.2908296e-33
+PUA = 3.1106794e-40
+UB = 1e-19
+UC = -2.3503344e-27
+LUC = 1.6694128e-34
+WUC = -1.3815828e-33
+PUC = 2.7982271e-40
+EU = 2.9
+VSAT = '103565.83*dvsatfactorn_hp'
+LVSAT = '-0.0022077023*dvsatfactorn_hp'
+WVSAT = '-0.00014346525*dvsatfactorn_hp'
+PVSAT = '5.9768831e-11*dvsatfactorn_hp'
+A0 = 0.98776623
+LA0 = 2.0797175e-07
+WA0 = 1.3811954e-06
+PA0 = -3.5288469e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8214409
+LPCLM = -1.0358339e-08
+WPCLM = -6.6575108e-10
+PPCLM = 2.7859261e-16
+PDIBLC1 = 0
+PDIBLC2 = 0.0057171013
+LPDIBLC2 = 1.1038475e-09
+WPDIBLC2 = 7.1689562e-11
+PPDIBLC2 = -2.98737e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72704928
+LPVAG = -2.0675964e-08
+WPVAG = -1.342734e-09
+PPVAG = 5.5954255e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7131625e-10
+LALPHA0 = -4.4153974e-17
+WALPHA0 = -2.8684438e-18
+PALPHA0 = 1.1951623e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165762
+LAIGC = 8.8245096e-12
+WAIGC = 5.6040334e-13
+PAIGC = -2.3573221e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5655024
+LUTE = 2.6933773e-08
+WUTE = 1.7481238e-09
+PUTE = -7.2862684e-16
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.315 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.38218008+dvth0n315_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-3.4809123e-09+dlvth0n315_hp'
+WVTH0 = '-3.9127609e-08+dwvth0n315_hp'
+PVTH0 = '4.310051e-15+dpvth0n315_hp'
+K1 = '0.7421651*dk1factorn_hp'
+LK1 = '-1.4410232e-08*dk1factorn_hp'
+WK1 = '-3.8951322e-08*dk1factorn_hp'
+PK1 = '6.2252204e-15*dk1factorn_hp'
+K2 = '-0.21194769*dk2factorn_hp'
+LK2 = '1.094607e-08*dk2factorn_hp'
+WK2 = '2.6429614e-08*dk2factorn_hp'
+PK2 = '-5.1963957e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.19411364
+LVOFF = 1.1762292e-08
+WVOFF = 3.932994e-08
+PVOFF = -6.9520839e-15
+NFACTOR = 0.4234354
+LNFACTOR = 1.2438682e-07
+WNFACTOR = 4.7274763e-07
+PNFACTOR = -7.5811273e-14
+ETA0 = 0
+ETAB = -0.073178918
+LETAB = -1.7299335e-13
+WETAB = -2.420241e-15
+U0 = '(0.034168398*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.6301417e-10*du0factorn_hp'
+WU0 = '-1.3820356e-09*du0factorn_hp'
+PU0 = '3.1091846e-16*du0factorn_hp'
+UA = 5.5042818e-28
+LUA = 2.3768403e-34
+WUA = 2.8291883e-33
+PUA = -4.5626706e-40
+UB = 1e-19
+UC = -4.7603239e-27
+LUC = 6.1395114e-34
+WUC = 8.5970749e-34
+PUC = -1.3589646e-40
+EU = 2.9
+VSAT = '68326.339*dvsatfactorn_hp'
+LVSAT = '0.0035106215*dvsatfactorn_hp'
+WVSAT = '0.032629259*dvsatfactorn_hp'
+PVSAT = '-5.2582723e-09*dvsatfactorn_hp'
+A0 = 2.469269
+LA0 = -1.6995575e-07
+WA0 = 3.3978703e-09
+PA0 = -1.4121123e-15
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8205068
+LPCLM = -9.968737e-09
+WPCLM = 2.0293963e-10
+PPCLM = -8.3737118e-17
+PDIBLC1 = 0
+PDIBLC2 = 0.0058169879
+LPDIBLC2 = 1.0622438e-09
+WPDIBLC2 = -2.1204921e-11
+PPDIBLC2 = 8.8177723e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72517829
+LPVAG = -1.9896681e-08
+WPVAG = 3.972899e-10
+PPVAG = -1.651905e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.6731878e-10
+LALPHA0 = -4.2489321e-17
+WALPHA0 = 8.4920858e-19
+PALPHA0 = -3.5296464e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010166516
+LAIGC = 8.5028221e-12
+WAIGC = -1.4120089e-13
+PAIGC = 6.3437211e-20
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7489339
+LUTE = 4.8834905e-08
+WUTE = 1.7233945e-07
+PUTE = -2.1096679e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.415 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.31924121+dvth0n415_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.4526445e-09+dlvth0n415_hp'
+WVTH0 = '-1.1938016e-08+dwvth0n415_hp'
+PVTH0 = '8.8275443e-16+dpvth0n415_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14614313*dk2factorn_hp'
+LK2 = '-7.4528309e-11*dk2factorn_hp'
+WK2 = '-1.9979575e-09*dk2factorn_hp'
+PK2 = '-4.3549727e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.095275885
+LVOFF = -7.4858222e-09
+WVOFF = -3.3679696e-09
+PVOFF = 1.3631012e-15
+NFACTOR = 1.8351123
+LNFACTOR = -1.1047043e-07
+WNFACTOR = -1.3709679e-07
+PNFACTOR = 2.5647061e-14
+ETA0 = 0
+ETAB = -0.073178568
+LETAB = -1.9503545e-13
+WETAB = -1.5361338e-13
+PETAB = 9.522188e-21
+U0 = '(0.032017379*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.2698238e-10*du0factorn_hp'
+WU0 = '-4.527954e-10*du0factorn_hp'
+PU0 = '1.6575273e-16*du0factorn_hp'
+UA = 9.7288564e-27
+LUA = -1.1588683e-33
+WUA = -1.1358927e-33
+PUA = 1.4704353e-40
+UB = 1e-19
+UC = -3.9124612e-27
+LUC = 4.1494924e-34
+WUC = 4.934308e-34
+PUC = -4.992764e-41
+EU = 2.9
+VSAT = '174591.49*dvsatfactorn_hp'
+LVSAT = '-0.014731039*dvsatfactorn_hp'
+WVSAT = '-0.013277285*dvsatfactorn_hp'
+PVSAT = '2.6221249e-09*dvsatfactorn_hp'
+A0 = 3.2319766
+LA0 = -2.946181e-07
+WA0 = -3.2609184e-07
+PA0 = 5.2442022e-14
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 2.0925426
+LPCLM = -7.7884726e-08
+WPCLM = -1.1731653e-07
+PPCLM = 2.925597e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.0063523223
+LPDIBLC2 = 9.5800059e-10
+WPDIBLC2 = -2.5246939e-10
+PPDIBLC2 = 5.385083e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 1.1674571
+LPVAG = -1.3048219e-07
+WPVAG = -1.9066716e-07
+PPVAG = 4.760775e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.019467252
+LPDITS = -2.3556416e-09
+WPDITS = -4.0898528e-09
+PPDITS = 1.0176372e-15
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.9881981e-11
+LALPHA0 = 6.7683549e-17
+WALPHA0 = 1.941419e-16
+PALPHA0 = -4.7947644e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.01004784
+LAIGC = 3.8263231e-11
+WAIGC = 5.1126708e-11
+PAIGC = -1.279306e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.3026638
+LUTE = -1.1778197e-08
+WUTE = -2.0449245e-08
+PUTE = 5.0881811e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.515 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30707474+dvth0n515_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.8713125e-09+dlvth0n515_hp'
+WVTH0 = '-9.7723845e-09+dwvth0n515_hp'
+PVTH0 = '1.1642315e-15+dpvth0n515_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14391341*dk2factorn_hp'
+LK2 = '-4.4448453e-09*dk2factorn_hp'
+WK2 = '-2.3948468e-09*dk2factorn_hp'
+PK2 = '3.4241915e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.14912264
+LVOFF = 7.2942693e-09
+WVOFF = 6.2167521e-09
+PVOFF = -1.2677551e-15
+NFACTOR = 1.0649056
+LNFACTOR = 3.361418e-08
+ETA0 = 0
+ETAB = -0.073179431
+LETAB = -1.4154001e-13
+U0 = '(0.030508025*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.0347498e-09*du0factorn_hp'
+WU0 = '-1.8413048e-10*du0factorn_hp'
+PU0 = '2.7393532e-16*du0factorn_hp'
+UA = 5.9720662e-27
+LUA = -9.8299338e-34
+WUA = -4.6718405e-34
+PUA = 1.157378e-40
+UB = 1e-19
+UC = -1.9877988e-27
+LUC = 2.8835331e-34
+WUC = 1.5084089e-34
+PUC = -2.7393564e-41
+EU = 2.9
+VSAT = '116067.3*dvsatfactorn_hp'
+LVSAT = '-0.015389625*dvsatfactorn_hp'
+WVSAT = '-0.0028599795*dvsatfactorn_hp'
+PVSAT = '2.7393532e-09*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.02196635
+LKETA = 7.6948124e-09
+WKETA = 1.4299897e-09
+PKETA = -1.3696766e-15
+DWG = 0
+DWB = 0
+PCLM = 1.433461
+LPCLM = 8.6474657e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0049339549
+LPDIBLC2 = 1.2605333e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.096293299
+LPVAG = 1.3697708e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0035094493
+LPDITS = 3.3614212e-09
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1105668e-09
+LALPHA0 = -2.0168524e-16
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010335069
+LAIGC = -3.360789e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4948602
+LUTE = 3.6044121e-08
+WUTE = 1.3761721e-08
+PUTE = -3.4241915e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.615 NMOS
+LMIN = '2.91000000e-07+dlminn_hp'
+LMAX = '2.95000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.27309323+dvth0n615_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.4548313e-08+dlvth0n615_hp'
+WVTH0 = '-6.5441407e-09+dwvth0n615_hp'
+PVTH0 = '-1.8450835e-15+dpvth0n615_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13866483*dk2factorn_hp'
+LK2 = '-3.1936459e-09*dk2factorn_hp'
+WK2 = '-2.8934616e-09*dk2factorn_hp'
+PK2 = '2.2355522e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.13116286
+LVOFF = -1.0055959e-08
+WVOFF = 4.5105729e-09
+PVOFF = 3.8051658e-16
+NFACTOR = 2.176957
+LNFACTOR = -1.074685e-07
+WNFACTOR = -1.0564488e-07
+PNFACTOR = 1.3402855e-14
+ETA0 = 0
+ETAB = -0.073177838
+LETAB = -5.3785205e-13
+WETAB = -1.5131277e-13
+PETAB = 3.7649643e-20
+U0 = '(-0.029989369*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.0553377e-08*du0factorn_hp'
+WU0 = '5.563122e-09*du0factorn_hp'
+PU0 = '-8.2693677e-16*du0factorn_hp'
+UA = -1.0786988e-26
+LUA = 8.8237554e-34
+WUA = 1.1249261e-33
+PUA = -6.1472246e-41
+UB = 1e-19
+UC = -4e-28
+EU = 2.9
+VSAT = '-84085.984*dvsatfactorn_hp'
+LVSAT = '0.045213605*dvsatfactorn_hp'
+WVSAT = '0.016154582*dvsatfactorn_hp'
+PVSAT = '-3.0179536e-09*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = -0.026874382
+LKETA = 9.7332682e-09
+WKETA = 6.0698593e-09
+PKETA = -1.5633299e-15
+DWG = 0
+DWB = 0
+PCLM = 0.35238129
+LPCLM = 3.5590079e-07
+WPCLM = 1.0270257e-07
+PPCLM = -2.5595483e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.00237793
+LPDIBLC2 = 1.8500079e-09
+WPDIBLC2 = 2.4282237e-10
+PPDIBLC2 = -5.600008e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = -1.6628168
+LPVAG = 5.7554963e-07
+WPVAG = 1.6711546e-07
+PPVAG = -4.1664392e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.041335907
+LPDITS = 1.2773401e-08
+WPDITS = 3.5935135e-09
+PPDITS = -8.9413804e-16
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 2.9149997e-09
+LALPHA0 = -6.488036e-16
+WALPHA0 = -1.7142112e-16
+PALPHA0 = 4.2476244e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010806271
+LAIGC = -1.512245e-10
+WAIGC = -4.4764224e-11
+PAIGC = 1.1173578e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.49
+WUTE = 1.33e-08
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.016 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.32499741+dvth0n016_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.6413937e-09+dlvth0n016_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.1140687
+LVOFF = 1.6657595e-09
+NFACTOR = 1.3186953
+LNFACTOR = -1.7855539e-10
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.032*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 4.1726935e-27
+LUA = -3.4996694e-34
+UB = 1e-19
+UC = -6.653969e-28
+LUC = -3.9371301e-35
+EU = 2.9
+VSAT = '90000*dvsatfactorn_hp'
+A0 = 1.7296625
+LA0 = 4.374607e-08
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8212218
+LPCLM = -1.0265312e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0057415631
+LPDIBLC2 = 1.0936518e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72659118
+LPVAG = -2.048501e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7033684e-10
+LALPHA0 = -4.3745908e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165933
+LAIGC = 8.7492141e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.461
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n016_hp'
+PVTH0 = '0.0+dpvth0n016_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.116 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.31634803+dvth0n116_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.4315591e-09+dlvth0n116_hp'
+WVTH0 = '8.5871027e-08+dwvth0n116_hp'
+PVTH0 = '-7.8447628e-15+dpvth0n116_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13507936*dk2factorn_hp'
+LK2 = '-4.5764656e-10*dk2factorn_hp'
+WK2 = '-4.8852081e-08*dk2factorn_hp'
+PK2 = '4.5435151e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10831835
+LVOFF = 2.0609101e-09
+WVOFF = -5.7089477e-08
+PVOFF = -3.9230558e-15
+NFACTOR = 1.3189862
+LNFACTOR = -2.5327874e-10
+WNFACTOR = -2.8886124e-09
+PNFACTOR = 7.4185343e-16
+ETA0 = 0
+ETAB = -0.073179891
+LETAB = 7.4723351e-14
+WETAB = 2.8886124e-12
+PETAB = -7.4185343e-19
+U0 = '(0.032365638*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0137943e-10*du0factorn_hp'
+WU0 = '-3.630058e-09*du0factorn_hp'
+PU0 = '1.999295e-15*du0factorn_hp'
+UA = 3.7119326e-27
+LUA = -2.9504528e-34
+WUA = 4.574434e-33
+PUA = -5.4526227e-40
+UB = 1e-19
+UC = 2.3712413e-28
+LUC = -1.6569038e-34
+WUC = -8.9602289e-33
+PUC = 1.2540958e-39
+EU = 2.9
+VSAT = '84343.372*dvsatfactorn_hp'
+LVSAT = '0.00091535426*dvsatfactorn_hp'
+WVSAT = '0.056159001*dvsatfactorn_hp'
+PVSAT = '-9.0876371e-09*dvsatfactorn_hp'
+A0 = 1.8427956
+LA0 = 2.5438849e-08
+WA0 = -1.1231853e-06
+PA0 = 1.8175409e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.8212218
+LPCLM = -1.0265312e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0057415631
+LPDIBLC2 = 1.0936518e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.72659118
+LPVAG = -2.048501e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.7033684e-10
+LALPHA0 = -4.3745908e-17
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010165933
+LAIGC = 8.7492141e-12
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4175179
+LUTE = -1.1167065e-08
+WUTE = -4.3168999e-07
+PUTE = 1.1086662e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.216 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.36144464+dvth0n216_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-1.3032636e-09+dlvth0n216_hp'
+WVTH0 = '-4.6216943e-08+dwvth0n216_hp'
+PVTH0 = '8.952533e-15+dpvth0n216_hp'
+K1 = '0.64228676*dk1factorn_hp'
+LK1 = '3.6671537e-10*dk1factorn_hp'
+WK1 = '2.8450081e-08*dk1factorn_hp'
+PK1 = '-1.0741093e-15*dk1factorn_hp'
+K2 = '-0.14789067*dk2factorn_hp'
+LK2 = '1.8684607e-09*dk2factorn_hp'
+WK2 = '-1.1327757e-08*dk2factorn_hp'
+PK2 = '-2.2696531e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.12688974
+LVOFF = 1.6547774e-09
+WVOFF = -2.693877e-09
+PVOFF = -2.7334932e-15
+NFACTOR = 1.4585529
+LNFACTOR = -1.0049934e-08
+WNFACTOR = -4.1167951e-07
+PNFACTOR = 2.9436258e-14
+ETA0 = 0
+ETAB = -0.073178728
+LETAB = -2.2386618e-13
+WETAB = -5.1676395e-13
+PETAB = 1.3271532e-19
+U0 = '(0.031427596*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '6.4532247e-10*du0factorn_hp'
+WU0 = '-8.8253077e-10*du0factorn_hp'
+PU0 = '-4.8069488e-16*du0factorn_hp'
+UA = 6.1599405e-27
+LUA = -6.1373016e-34
+WUA = -2.595781e-33
+PUA = 3.8816576e-40
+UB = 1e-19
+UC = -2.9044764e-27
+LUC = 3.0703948e-34
+WUC = 2.4151918e-34
+PUC = -1.3052994e-40
+EU = 2.9
+VSAT = '107107.12*dvsatfactorn_hp'
+LVSAT = '-0.0031030109*dvsatfactorn_hp'
+WVSAT = '-0.010516006*dvsatfactorn_hp'
+PVSAT = '2.6821545e-09*dvsatfactorn_hp'
+A0 = 1.0809095
+LA0 = 1.8442326e-07
+WA0 = 1.108379e-06
+PA0 = -2.8391125e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.9122459
+LPCLM = -3.3315668e-08
+WPCLM = -2.6660951e-07
+PPCLM = 6.7514494e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.0059272359
+LPDIBLC2 = 1.0507213e-09
+WPDIBLC2 = -5.4383548e-10
+PPDIBLC2 = 1.2574334e-16
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.87453352
+LPVAG = -5.7962928e-08
+WPVAG = -4.3332311e-07
+PPVAG = 1.0977282e-13
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.013169339
+LPDITS = -8.0127232e-10
+WPDITS = -9.2829944e-09
+PPDITS = 2.3469266e-15
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 3.2028936e-10
+LALPHA0 = -5.9713555e-18
+WALPHA0 = 4.3948907e-16
+PALPHA0 = -1.1064166e-22
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010126213
+LAIGC = 1.8823314e-11
+WAIGC = 1.1633964e-10
+PAIGC = -2.9507039e-17
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5611641
+LUTE = 2.5836979e-08
+WUTE = -1.0950252e-08
+PUTE = 2.4817765e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.316 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.33318314+dvth0n316_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '8.9064934e-09+dlvth0n316_hp'
+WVTH0 = '-1.9933747e-08+dwvth0n316_hp'
+PVTH0 = '-5.42541e-16+dpvth0n316_hp'
+K1 = '0.69098949*dk1factorn_hp'
+LK1 = '-1.4720161e-09*dk1factorn_hp'
+WK1 = '-1.6843461e-08*dk1factorn_hp'
+PK1 = '6.3591096e-16*dk1factorn_hp'
+K2 = '-0.16944301*dk2factorn_hp'
+LK2 = '2.000368e-10*dk2factorn_hp'
+WK2 = '8.7159171e-09*dk2factorn_hp'
+PK2 = '-7.180189e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.1492897
+LVOFF = 4.2990388e-10
+WVOFF = 1.8138092e-08
+PVOFF = -1.5943608e-15
+NFACTOR = 0.68835983
+LNFACTOR = 5.7408628e-08
+WNFACTOR = 3.0460007e-07
+PNFACTOR = -3.3300205e-14
+ETA0 = 0
+ETAB = -0.073179448
+LETAB = -3.8918425e-14
+WETAB = 1.5297133e-13
+PETAB = -3.9286097e-20
+U0 = '(0.030918248*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '5.868879e-11*du0factorn_hp'
+WU0 = '-4.0883724e-10*du0factorn_hp'
+PU0 = '6.4874442e-17*du0factorn_hp'
+UA = 1.0926856e-27
+LUA = 1.005905e-34
+WUA = 2.116766e-33
+PUA = -2.7615245e-40
+UB = 1e-19
+UC = -2.9080765e-27
+LUC = 1.4566594e-34
+WUC = 2.4486723e-34
+PUC = 1.9547452e-41
+EU = 2.9
+VSAT = '67371.516*dvsatfactorn_hp'
+LVSAT = '0.0037520198*dvsatfactorn_hp'
+WVSAT = '0.026438102*dvsatfactorn_hp'
+PVSAT = '-3.6930241e-09*dvsatfactorn_hp'
+A0 = 2.1830575
+LA0 = -9.7595775e-08
+WA0 = 8.3381383e-08
+PA0 = -2.1633544e-14
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.5408765
+LPCLM = 6.0727392e-08
+WPCLM = 7.8764028e-08
+PPCLM = -1.9945551e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.0051652384
+LPDIBLC2 = 1.2270191e-09
+WPDIBLC2 = 1.6482213e-10
+PPDIBLC2 = -3.8213587e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.27094696
+LPVAG = 9.4942084e-08
+WPVAG = 1.2801239e-07
+PPVAG = -3.242884e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.00023706745
+LPDITS = 2.4682646e-09
+WPDITS = 2.7440183e-09
+PPDITS = -6.9374271e-16
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 9.3272284e-10
+LALPHA0 = -1.6015278e-16
+WALPHA0 = -1.3007406e-16
+PALPHA0 = 3.2747057e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010288284
+LAIGC = -2.2282656e-11
+WAIGC = -3.4387211e-11
+PAIGC = 8.7215135e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7219471
+LUTE = 4.2012088e-08
+WUTE = 1.3857786e-07
+PUTE = -1.2561075e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.416 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.31147433+dvth0n416_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '6.4162671e-09+dlvth0n416_hp'
+WVTH0 = '-1.055554e-08+dwvth0n416_hp'
+PVTH0 = '5.3323675e-16+dpvth0n416_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14359038*dk2factorn_hp'
+LK2 = '-7.1991309e-10*dk2factorn_hp'
+WK2 = '-2.452418e-09*dk2factorn_hp'
+PK2 = '-3.2060055e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.10247279
+LVOFF = -5.6663013e-09
+WVOFF = -2.0868156e-09
+PVOFF = 1.0391998e-15
+NFACTOR = 1.6236933
+LNFACTOR = -5.7019472e-08
+WNFACTOR = -9.9463975e-08
+PNFACTOR = 1.6132734e-14
+ETA0 = 0
+ETAB = -0.073178826
+LETAB = -1.2985846e-13
+WETAB = -1.1594948e-13
+U0 = '(0.030321041*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.8857596e-12*du0factorn_hp'
+WU0 = '-1.5084391e-10*du0factorn_hp'
+PU0 = '8.9413351e-17*du0factorn_hp'
+UA = 7.8463111e-27
+LUA = -6.8292317e-34
+WUA = -8.0080023e-34
+PUA = 6.2325454e-41
+UB = 1e-19
+UC = -3.1828134e-27
+LUC = 2.3047966e-34
+WUC = 3.6355357e-34
+PUC = -1.7092078e-41
+EU = 2.9
+VSAT = '148592.9*dvsatfactorn_hp'
+LVSAT = '-0.0081580769*dvsatfactorn_hp'
+WVSAT = '-0.0086495368*dvsatfactorn_hp'
+PVSAT = '1.4521377e-09*dvsatfactorn_hp'
+A0 = 3.0600875
+LA0 = -2.511611e-07
+WA0 = -2.9549558e-07
+PA0 = 4.4706675e-14
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.9262413
+LPCLM = -3.5840425e-08
+WPCLM = -8.7713551e-08
+PPCLM = 2.1771745e-14
+PDIBLC1 = 0
+PDIBLC2 = 0.0059762238
+LPDIBLC2 = 1.0530858e-09
+WPDIBLC2 = -1.8552353e-10
+PPDIBLC2 = 3.6925576e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.89732801
+LPVAG = -6.2188154e-08
+WPVAG = -1.4258422e-07
+PPVAG = 3.5451423e-14
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0.013665803
+LPDITS = -8.8891941e-10
+WPDITS = -3.0571956e-09
+PPDITS = 7.5656078e-16
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 2.9598925e-10
+LALPHA0 = -2.1218911e-18
+WALPHA0 = 1.4499485e-16
+PALPHA0 = -3.5522285e-23
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.01012009
+LAIGC = 1.9997053e-11
+WAIGC = 3.8272747e-11
+PAIGC = -9.5433211e-18
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.389685
+LUTE = 1.0222494e-08
+WUTE = -4.9593659e-09
+PUTE = 1.1720299e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.516 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30707449+dvth0n516_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.871376e-09+dlvth0n516_hp'
+WVTH0 = '-9.7723681e-09+dwvth0n516_hp'
+PVTH0 = '1.1642274e-15+dpvth0n516_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14391389*dk2factorn_hp'
+LK2 = '-4.4447247e-09*dk2factorn_hp'
+WK2 = '-2.3948341e-09*dk2factorn_hp'
+PK2 = '3.4241592e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.14912169
+LVOFF = 7.2940307e-09
+WVOFF = 6.2166895e-09
+PVOFF = -1.2677392e-15
+NFACTOR = 1.0649069
+LNFACTOR = 3.3613864e-08
+ETA0 = 0
+ETAB = -0.073179477
+LETAB = -1.2985846e-13
+U0 = '(0.03050806*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.0347586e-09*du0factorn_hp'
+WU0 = '-1.8413335e-10*du0factorn_hp'
+PU0 = '2.7393605e-16*du0factorn_hp'
+UA = 5.9720637e-27
+LUA = -9.8299275e-34
+WUA = -4.671842e-34
+PUA = 1.1573784e-40
+UB = 1e-19
+UC = -1.9877977e-27
+LUC = 2.8835304e-34
+WUC = 1.5084079e-34
+PUC = -2.7393538e-41
+EU = 2.9
+VSAT = '116067.46*dvsatfactorn_hp'
+LVSAT = '-0.015389666*dvsatfactorn_hp'
+WVSAT = '-0.0028600082*dvsatfactorn_hp'
+PVSAT = '2.7393605e-09*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.021966269
+LKETA = 7.6948328e-09
+WKETA = 1.4300041e-09
+PKETA = -1.3696802e-15
+DWG = 0
+DWB = 0
+PCLM = 1.4334685
+LPCLM = 8.6472752e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0049339568
+LPDIBLC2 = 1.2605329e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.096293037
+LPVAG = 1.3697714e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0035094529
+LPDITS = 3.3614221e-09
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.110567e-09
+LALPHA0 = -2.0168529e-16
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010335106
+LAIGC = -3.361711e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4948589
+LUTE = 3.6043781e-08
+WUTE = 1.3761594e-08
+PUTE = -3.4241592e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.616 NMOS
+LMIN = '2.95000000e-07+dlminn_hp'
+LMAX = '2.99000000e-07+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.2394504+dvth0n616_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.3053892e-08+dlvth0n616_hp'
+WVTH0 = '-3.3480797e-09+dwvth0n616_hp'
+PVTH0 = '-2.6531117e-15+dpvth0n616_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.10062416*dk2factorn_hp'
+LK2 = '-1.2811089e-08*dk2factorn_hp'
+WK2 = '-6.5073583e-09*dk2factorn_hp'
+PK2 = '1.1372206e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.060974225
+LVOFF = -2.7801048e-08
+WVOFF = -2.1573199e-09
+PVOFF = 2.0662933e-15
+NFACTOR = 0.86622641
+LNFACTOR = 2.2391041e-07
+WNFACTOR = 1.8874646e-08
+PNFACTOR = -1.8078172e-14
+ETA0 = 0
+ETAB = -0.073179452
+LETAB = -1.2985846e-13
+WETAB = -2.394e-15
+U0 = '(0.013256952*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.8015741e-10*du0factorn_hp'
+WU0 = '1.454722e-09*du0factorn_hp'
+PU0 = '2.1174893e-16*du0factorn_hp'
+UA = -5.8881766e-27
+LUA = -3.5614203e-34
+WUA = 6.5953864e-34
+PUA = 5.6187021e-41
+UB = 1e-19
+UC = -1.5412323e-27
+LUC = 2.8852635e-34
+WUC = 1.0841707e-34
+PUC = -2.7410004e-41
+EU = 2.9
+VSAT = '-107343.97*dvsatfactorn_hp'
+LVSAT = '0.05109369*dvsatfactorn_hp'
+WVSAT = '0.018364078*dvsatfactorn_hp'
+PVSAT = '-3.5765583e-09*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.036589832
+LKETA = -6.3117544e-09
+WKETA = 4.0765624e-11
+PKETA = -3.9054446e-17
+DWG = 0
+DWB = 0
+PCLM = 1.4389981
+LPCLM = 8.1182318e-08
+WPCLM = -5.2531329e-10
+PPCLM = 5.0259122e-16
+PDIBLC1 = 0
+PDIBLC2 = 0.0050144442
+LPDIBLC2 = 1.1834443e-09
+WPDIBLC2 = -7.6463031e-12
+PPDIBLC2 = 7.3234103e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.10503778
+LPVAG = 1.2860062e-07
+WPVAG = -8.3075032e-10
+PPVAG = 7.9576943e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0032948436
+LPDITS = 3.1558587e-09
+WPDITS = -2.0387882e-11
+PPDITS = 1.9528518e-17
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.0976901e-09
+LALPHA0 = -1.893514e-16
+WALPHA0 = 1.2233076e-18
+PALPHA0 = -1.1717197e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010332999
+LAIGC = -3.1571839e-11
+WAIGC = 2.0009185e-13
+PAIGC = -1.9430073e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.2997991
+LUTE = -4.808659e-08
+WUTE = -4.7690847e-09
+PUTE = 4.568226e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.017 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.28794191+dvth0n017_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.3157989e-08+dlvth0n017_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13316819*dk2factorn_hp'
+LK2 = '-1.7545459e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.08815765
+LVOFF = -4.9887157e-09
+NFACTOR = 1.318
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.032*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 4.1626987e-27
+LUA = -3.4740008e-34
+UB = 1e-19
+UC = -1.8848725e-27
+LUC = 2.7381443e-34
+EU = 2.9
+VSAT = '90000*dvsatfactorn_hp'
+A0 = 2.0366362
+LA0 = -3.5090918e-08
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4294059
+LPCLM = 9.0360867e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0048761412
+LPDIBLC2 = 1.3159094e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.090000834
+LPVAG = 1.4300412e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0036636234
+LPDITS = 3.5090918e-09
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1198174e-09
+LALPHA0 = -2.1054551e-16
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010336636
+LAIGC = -3.5090918e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6509244
+LUTE = 4.8776375e-08
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n017_hp'
+PVTH0 = '0.0+dpvth0n017_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.117 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.28959044+dvth0n117_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.1303445e-08+dlvth0n117_hp'
+WVTH0 = '-1.6366624e-08+dwvth0n117_hp'
+PVTH0 = '1.8411911e-14+dpvth0n117_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13145904*dk2factorn_hp'
+LK2 = '-1.3874174e-09*dk2factorn_hp'
+WK2 = '-1.69684e-08*dk2factorn_hp'
+PK2 = '-3.6448518e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.083493581
+LVOFF = -4.3145861e-09
+WVOFF = -4.630487e-08
+PVOFF = -6.6927586e-15
+NFACTOR = 1.3854732
+LNFACTOR = -1.7328466e-08
+WNFACTOR = -6.6987387e-07
+PNFACTOR = 1.7203701e-13
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.033296932*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.4055421e-10*du0factorn_hp'
+WU0 = '-1.2875939e-08*du0factorn_hp'
+PU0 = '4.3738222e-15*du0factorn_hp'
+UA = 4.7106019e-27
+LUA = -5.5152354e-34
+WUA = -5.4395832e-33
+PUA = 2.0265376e-39
+UB = 1e-19
+UC = -2.0353239e-27
+LUC = 4.1791971e-34
+WUC = 1.4936807e-33
+PUC = -1.4306772e-39
+EU = 2.9
+VSAT = '90766.592*dvsatfactorn_hp'
+LVSAT = '-0.00073425702*dvsatfactorn_hp'
+WVSAT = '-0.007610724*dvsatfactorn_hp'
+PVSAT = '7.2897037e-09*dvsatfactorn_hp'
+A0 = 2.0213044
+LA0 = -2.0405777e-08
+WA0 = 1.5221448e-07
+PA0 = -1.4579407e-13
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4294059
+LPCLM = 9.0360867e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0048761412
+LPDIBLC2 = 1.3159094e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.090000834
+LPVAG = 1.4300412e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0036636234
+LPDITS = 3.5090918e-09
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1198174e-09
+LALPHA0 = -2.1054551e-16
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010336636
+LAIGC = -3.5090918e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6509244
+LUTE = 4.8776375e-08
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.217 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.284287+dvth0n217_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.8512362e-08+dlvth0n217_hp'
+WVTH0 = '-8.3286252e-10+dwvth0n217_hp'
+PVTH0 = '-2.7030066e-15+dpvth0n217_hp'
+K1 = '0.65503543*dk1factorn_hp'
+LK1 = '-2.9073991e-09*dk1factorn_hp'
+WK1 = '-8.8907854e-09*dk1factorn_hp'
+PK1 = '8.5157721e-15*dk1factorn_hp'
+K2 = '-0.13754971*dk2factorn_hp'
+LK2 = '-7.8730537e-10*dk2factorn_hp'
+WK2 = '8.7116384e-10*dk2factorn_hp'
+PK2 = '-5.4025799e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.095372489
+LVOFF = -6.439482e-09
+WVOFF = -1.1511549e-08
+PVOFF = -4.6893862e-16
+NFACTOR = 1.1831801
+LNFACTOR = 6.0671301e-08
+WNFACTOR = -7.7357537e-08
+PNFACTOR = -5.642431e-14
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.029192085*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.2194463e-09*du0factorn_hp'
+WU0 = '-8.5284256e-10*du0factorn_hp'
+PU0 = '-4.8831941e-16*du0factorn_hp'
+UA = 2.7178235e-27
+LUA = 2.7027432e-34
+WUA = 3.9726492e-34
+PUA = -3.8050829e-40
+UB = 1e-19
+UC = -1.5587247e-27
+LUC = -3.857648e-35
+WUC = 9.7721803e-35
+PUC = -9.3599897e-41
+EU = 2.9
+VSAT = '88159.146*dvsatfactorn_hp'
+LVSAT = '0.0017632069*dvsatfactorn_hp'
+WVSAT = '2.648513e-05*dvsatfactorn_hp'
+PVSAT = '-2.5367987e-11*dvsatfactorn_hp'
+A0 = 2.0736342
+LA0 = -7.0528277e-08
+WA0 = -1.0594152e-09
+PA0 = 1.0147291e-15
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4289402
+LPCLM = 9.0806911e-08
+WPCLM = 1.3639952e-09
+PPCLM = -1.3064619e-15
+PDIBLC1 = 0
+PDIBLC2 = 0.0048693595
+LPDIBLC2 = 1.3224051e-09
+WPDIBLC2 = 1.9863748e-11
+PPDIBLC2 = -1.9025895e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.089263839
+LPVAG = 1.4371003e-07
+WPVAG = 2.1586589e-09
+PPVAG = -2.0676067e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0036817081
+LPDITS = 3.5264136e-09
+WPDITS = 5.2970011e-11
+PPDITS = -5.0735736e-17
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1209025e-09
+LALPHA0 = -2.1158482e-16
+WALPHA0 = -3.1782006e-18
+PALPHA0 = 3.0441441e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010336817
+LAIGC = -3.5264131e-11
+WAIGC = -5.2968263e-13
+PAIGC = 5.0734062e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6828691
+LUTE = 5.7093256e-08
+WUTE = 9.356622e-08
+PUTE = -2.4360144e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.317 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29211192+dvth0n317_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.9454405e-08+dlvth0n317_hp'
+WVTH0 = '-8.1100351e-09+dwvth0n317_hp'
+PVTH0 = '-3.5791068e-15+dpvth0n317_hp'
+K1 = '0.6398156*dk1factorn_hp'
+LK1 = '1.1670464e-08*dk1factorn_hp'
+WK1 = '5.2636615e-09*dk1factorn_hp'
+PK1 = '-5.0416403e-15*dk1factorn_hp'
+K2 = '-0.1295397*dk2factorn_hp'
+LK2 = '-1.004793e-08*dk2factorn_hp'
+WK2 = '-6.5781406e-09*dk2factorn_hp'
+PK2 = '3.209801e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.097124426
+LVOFF = -1.2967183e-08
+WVOFF = -9.8822481e-09
+PVOFF = 5.6018228e-15
+NFACTOR = 1.1689141
+LNFACTOR = -6.6007325e-08
+WNFACTOR = -6.4090134e-08
+PNFACTOR = 6.1386812e-14
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.029398783*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '4.4891776e-10*du0factorn_hp'
+WU0 = '-1.0450717e-09*du0factorn_hp'
+PU0 = '2.2827217e-16*du0factorn_hp'
+UA = 3.5552724e-27
+LUA = -5.3185104e-34
+WUA = -3.8156261e-34
+PUA = 3.654683e-40
+UB = 1e-19
+UC = -1.800127e-27
+LUC = -1.3887765e-34
+WUC = 3.2222594e-34
+PUC = -3.1981233e-43
+EU = 2.9
+VSAT = '92937.842*dvsatfactorn_hp'
+LVSAT = '-0.002813924*dvsatfactorn_hp'
+WVSAT = '-0.0044177024*dvsatfactorn_hp'
+PVSAT = '4.2313637e-09*dvsatfactorn_hp'
+A0 = 2.0721583
+LA0 = -6.9114625e-08
+WA0 = 3.1317719e-10
+PA0 = -2.9996738e-16
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4308404
+LPCLM = 8.8986877e-08
+WPCLM = -4.0317573e-10
+PPCLM = 3.8616978e-16
+PDIBLC1 = 0
+PDIBLC2 = 0.004897032
+LPDIBLC2 = 1.2958999e-09
+WPDIBLC2 = -5.8716586e-12
+PPDIBLC2 = 5.623992e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.092271097
+LPVAG = 1.4082962e-07
+WPVAG = -6.3809114e-10
+PPVAG = 6.1117646e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0036079148
+LPDITS = 3.4557329e-09
+WPDITS = -1.5657736e-11
+PPDITS = 1.4997293e-17
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1164749e-09
+LALPHA0 = -2.0734398e-16
+WALPHA0 = 9.394636e-19
+PALPHA0 = -8.9983702e-25
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010336079
+LAIGC = -3.4557269e-11
+WAIGC = 1.5664771e-13
+PAIGC = -1.5004031e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6062006
+LUTE = 1.2286093e-08
+WUTE = 2.2264519e-08
+PUTE = 1.7310518e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.417 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.28817096+dvth0n417_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.2401038e-08+dlvth0n417_hp'
+WVTH0 = '-6.4075412e-09+dwvth0n417_hp'
+PVTH0 = '-5.3205218e-16+dpvth0n417_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13593624*dk2factorn_hp'
+LK2 = '-2.6856504e-09*dk2factorn_hp'
+WK2 = '-3.8148383e-09*dk2factorn_hp'
+PK2 = '2.9296233e-17*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.12406675
+LVOFF = -1.2053904e-10
+WVOFF = 1.7568375e-09
+PVOFF = 5.2072866e-17
+NFACTOR = 0.9894787
+LNFACTOR = 1.0585951e-07
+WNFACTOR = 1.3425969e-08
+PNFACTOR = -1.2859662e-14
+ETA0 = 0
+ETAB = -0.073179698
+LETAB = 9.4184575e-14
+WETAB = 4.2479523e-14
+PETAB = -4.0687737e-20
+U0 = '(0.025231909*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.3088767e-09*du0factorn_hp'
+WU0 = '7.5501788e-10*du0factorn_hp'
+PU0 = '-1.4323008e-16*du0factorn_hp'
+UA = 2.1987069e-27
+LUA = 7.6749454e-34
+WUA = 2.044737e-34
+PUA = -1.95849e-40
+UB = 1e-19
+UC = -9.9386473e-28
+LUC = -3.3168613e-34
+WUC = -2.6079363e-35
+PUC = 8.2973451e-41
+EU = 2.9
+VSAT = '70596.242*dvsatfactorn_hp'
+LVSAT = '0.011873026*dvsatfactorn_hp'
+WVSAT = '0.005233869*dvsatfactorn_hp'
+PVSAT = '-2.1133986e-09*dvsatfactorn_hp'
+A0 = 2.5444313
+LA0 = -1.1873026e-07
+WA0 = -2.0370877e-07
+PA0 = 2.1133986e-14
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4274145
+LPCLM = 9.2268281e-08
+WPCLM = 1.0768171e-09
+PPCLM = -1.0313969e-15
+PDIBLC1 = 0
+PDIBLC2 = 0.0048480391
+LPDIBLC2 = 1.3428262e-09
+WPDIBLC2 = 1.529326e-11
+PPDIBLC2 = -1.4648191e-17
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.086940222
+LPVAG = 1.4593564e-07
+WPVAG = 1.6648468e-09
+PPVAG = -1.5946236e-15
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0037385624
+LPDITS = 3.5808698e-09
+WPDITS = 4.0782017e-11
+PPDITS = -3.9061831e-17
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1243137e-09
+LALPHA0 = -2.1485219e-16
+WALPHA0 = -2.4469203e-18
+PALPHA0 = 2.3437092e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010337386
+LAIGC = -3.5808806e-11
+WAIGC = -4.078256e-13
+PAIGC = 3.9062352e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.650751
+LUTE = 7.7269467e-08
+WUTE = 4.151026e-08
+PUTE = -1.0762299e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.517 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.30707446+dvth0n517_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.8713845e-09+dlvth0n517_hp'
+WVTH0 = '-9.7723632e-09+dwvth0n517_hp'
+PVTH0 = '1.1642261e-15+dpvth0n517_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14391371*dk2factorn_hp'
+LK2 = '-4.4447703e-09*dk2factorn_hp'
+WK2 = '-2.3948483e-09*dk2factorn_hp'
+PK2 = '3.4241957e-16*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.14912242
+LVOFF = 7.2942165e-09
+WVOFF = 6.2167455e-09
+PVOFF = -1.2677536e-15
+NFACTOR = 1.0649055
+LNFACTOR = 3.3614222e-08
+ETA0 = 0
+ETAB = -0.07317946
+LETAB = -1.3439821e-13
+U0 = '(0.030508029*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.0347506e-09*du0factorn_hp'
+WU0 = '-1.8413155e-10*du0factorn_hp'
+PU0 = '2.7393559e-16*du0factorn_hp'
+UA = 5.9720647e-27
+LUA = -9.8299299e-34
+WUA = -4.6718399e-34
+PUA = 1.1573778e-40
+UB = 1e-19
+UC = -1.9877986e-27
+LUC = 2.8835325e-34
+WUC = 1.5084087e-34
+PUC = -2.7393559e-41
+EU = 2.9
+VSAT = '116067.36*dvsatfactorn_hp'
+LVSAT = '-0.01538964*dvsatfactorn_hp'
+WVSAT = '-0.0028599902*dvsatfactorn_hp'
+PVSAT = '2.7393559e-09*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.02196632
+LKETA = 7.6948198e-09
+WKETA = 1.4299951e-09
+PKETA = -1.3696779e-15
+DWG = 0
+DWB = 0
+PCLM = 1.433464
+LPCLM = 8.6473917e-08
+PDIBLC1 = 0
+PDIBLC2 = 0.0049339563
+LPDIBLC2 = 1.260533e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.096293294
+LPVAG = 1.3697708e-07
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0035094499
+LPDITS = 3.3614213e-09
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.110567e-09
+LALPHA0 = -2.0168528e-16
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010335095
+LAIGC = -3.3614292e-11
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.4948604
+LUTE = 3.6044165e-08
+WUTE = 1.3761736e-08
+PUTE = -3.4241957e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.617 NMOS
+LMIN = '2.99000000e-07+dlminn_hp'
+LMAX = '1.00000000e-06+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.23945002+dvth0n617_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.305399e-08+dlvth0n617_hp'
+WVTH0 = '-3.3480417e-09+dwvth0n617_hp'
+PVTH0 = '-2.6531214e-15+dpvth0n617_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.10062496*dk2factorn_hp'
+LK2 = '-1.2810885e-08*dk2factorn_hp'
+WK2 = '-6.5072799e-09*dk2factorn_hp'
+PK2 = '1.1372004e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.060974824
+LVOFF = -2.7800894e-08
+WVOFF = -2.1572758e-09
+PVOFF = 2.0662819e-15
+NFACTOR = 0.86623014
+LNFACTOR = 2.2390945e-07
+WNFACTOR = 1.8874158e-08
+PNFACTOR = -1.8078046e-14
+ETA0 = 0
+ETAB = -0.073179469
+LETAB = -1.255553e-13
+WETAB = 8.7707144e-16
+PETAB = -8.4007657e-22
+U0 = '(0.013256879*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.8013879e-10*du0factorn_hp'
+WU0 = '1.4547277e-09*du0factorn_hp'
+PU0 = '2.1174746e-16*du0factorn_hp'
+UA = -5.8881735e-27
+LUA = -3.5614282e-34
+WUA = 6.5953865e-34
+PUA = 5.6187018e-41
+UB = 1e-19
+UC = -1.5412323e-27
+LUC = 2.8852636e-34
+WUC = 1.0841707e-34
+PUC = -2.7410004e-41
+EU = 2.9
+VSAT = '-107343.64*dvsatfactorn_hp'
+LVSAT = '0.051093604*dvsatfactorn_hp'
+WVSAT = '0.018364055*dvsatfactorn_hp'
+PVSAT = '-3.5765522e-09*dvsatfactorn_hp'
+A0 = 1.4
+AGS = 0.6
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.036589663
+LKETA = -6.3117111e-09
+WKETA = 4.0777488e-11
+PKETA = -3.9057493e-17
+DWG = 0
+DWB = 0
+PCLM = 1.4389851
+LPCLM = 8.1185659e-08
+WPCLM = -5.2450821e-10
+PPCLM = 5.0238446e-16
+PDIBLC1 = 0
+PDIBLC2 = 0.0050144381
+LPDIBLC2 = 1.1834459e-09
+WPDIBLC2 = -7.6457728e-12
+PPDIBLC2 = 7.3232741e-18
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.10503894
+LPVAG = 1.2860033e-07
+WPVAG = -8.3083613e-10
+PPVAG = 7.9579146e-16
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = -0.0032948317
+LPDITS = 3.1558557e-09
+WPDITS = -2.0388734e-11
+PPDITS = 1.9528737e-17
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.0976899e-09
+LALPHA0 = -1.8935135e-16
+WALPHA0 = 1.2233237e-18
+PALPHA0 = -1.1717239e-24
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010332949
+LAIGC = -3.1558806e-11
+WAIGC = 2.0387038e-13
+PAIGC = -1.9527113e-19
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.2997946
+LUTE = -4.8087751e-08
+WUTE = -4.7695145e-09
+PUTE = 4.5683364e-15
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.018 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.262223+dvth0n018_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.7792074e-08+dlvth0n018_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.079550691
+LVOFF = -1.3232633e-08
+NFACTOR = 1.1434886
+LNFACTOR = 1.6715049e-07
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.032*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 2.616872e-27
+LUA = 1.1332237e-33
+UB = 1e-19
+UC = -1.4525879e-27
+LUC = -1.4023643e-34
+EU = 2.9
+VSAT = '104789.1*dvsatfactorn_hp'
+LVSAT = '-0.014165296*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.747891
+LUTE = 1.4165296e-07
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n018_hp'
+PVTH0 = '0.0+dpvth0n018_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.118 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.25890176+dvth0n118_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.0697671e-08+dlvth0n118_hp'
+WVTH0 = '3.2973208e-08+dwvth0n118_hp'
+PVTH0 = '-2.8846767e-14+dpvth0n118_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13600209*dk2factorn_hp'
+LK2 = '2.9640057e-09*dk2factorn_hp'
+WK2 = '9.9487623e-09*dk2factorn_hp'
+PK2 = '-2.9426648e-14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.075328597
+LVOFF = -1.2135172e-08
+WVOFF = -4.1916953e-08
+PVOFF = -1.0895593e-14
+NFACTOR = 1.1198393
+LNFACTOR = 2.3710102e-07
+WNFACTOR = 2.3479079e-07
+PNFACTOR = -6.944689e-13
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.031599163*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.1856023e-09*du0factorn_hp'
+WU0 = '3.9795049e-09*du0factorn_hp'
+PU0 = '-1.1770659e-14*du0factorn_hp'
+UA = 2.1470841e-27
+LUA = 1.9038651e-33
+WUA = 4.6640544e-33
+PUA = -7.6509285e-39
+UB = 1e-19
+UC = -1.4525879e-27
+LUC = -1.4023643e-34
+EU = 2.9
+VSAT = '104789.1*dvsatfactorn_hp'
+LVSAT = '-0.014165296*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7788363
+LUTE = 1.7129301e-07
+WUTE = 3.0722524e-07
+PUTE = -2.9426648e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.218 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26652666+dvth0n218_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.5523574e-08+dlvth0n218_hp'
+WVTH0 = '1.0639887e-08+dwvth0n218_hp'
+PVTH0 = '-1.3691835e-14+dpvth0n218_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12994508*dk2factorn_hp'
+LK2 = '-8.0711715e-09*dk2factorn_hp'
+WK2 = '-7.7922235e-09*dk2factorn_hp'
+PK2 = '2.8953857e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.077841127
+LVOFF = -2.3231371e-08
+WVOFF = -3.4557752e-08
+PVOFF = 2.1605175e-14
+NFACTOR = 1.1777195
+LNFACTOR = 6.5901576e-08
+WNFACTOR = 6.5259453e-08
+PNFACTOR = -1.9302572e-13
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.033423053*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.8330592e-09*du0factorn_hp'
+WU0 = '-1.3626663e-09*du0factorn_hp'
+PU0 = '6.6969248e-30*du0factorn_hp'
+UA = 3.739455e-27
+LUA = -7.0826479e-34
+UB = 1e-19
+UC = -1.1085693e-27
+LUC = -4.6974431e-34
+WUC = -1.0076304e-33
+PUC = 9.6512858e-40
+EU = 2.9
+VSAT = '104789.1*dvsatfactorn_hp'
+LVSAT = '-0.014165296*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6972071
+LUTE = 7.0826479e-08
+WUTE = 6.8133317e-08
+PUTE = 4.2860319e-28
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.318 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29111048+dvth0n318_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0413608e-08+dlvth0n318_hp'
+WVTH0 = '-1.2223063e-08+dwvth0n318_hp'
+PVTH0 = '3.6043312e-16+dpvth0n318_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13036375*dk2factorn_hp'
+LK2 = '-9.2586421e-09*dk2factorn_hp'
+WK2 = '-7.4028596e-09*dk2factorn_hp'
+PK2 = '3.9997334e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11260639
+LVOFF = 1.8617499e-09
+WVOFF = -2.2260598e-09
+PVOFF = -1.7314274e-15
+NFACTOR = 1.247891
+LNFACTOR = -1.4165296e-07
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.0341082*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.0618559e-09*du0factorn_hp'
+WU0 = '-1.9998532e-09*du0factorn_hp'
+PU0 = '1.142781e-15*du0factorn_hp'
+UA = 4.252619e-27
+LUA = -1.1997835e-33
+WUA = -4.7724248e-34
+PUA = 4.5711239e-40
+UB = 1e-19
+UC = -2.0262824e-27
+LUC = 7.773846e-35
+WUC = -1.5415732e-34
+PUC = 4.5596961e-40
+EU = 2.9
+VSAT = '104789.1*dvsatfactorn_hp'
+LVSAT = '-0.014165296*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7314645
+LUTE = 1.3226632e-07
+WUTE = 9.9992659e-08
+PUTE = -5.7139048e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.418 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.3069173+dvth0n418_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-5.5545805e-09+dlvth0n418_hp'
+WVTH0 = '-1.9051611e-08+dwvth0n418_hp'
+PVTH0 = '1.157869e-14+dpvth0n418_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14392216*dk2factorn_hp'
+LK2 = '4.9634304e-09*dk2factorn_hp'
+WK2 = '-1.5456247e-09*dk2factorn_hp'
+PK2 = '-2.1442019e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.14526691
+LVOFF = 2.0185391e-08
+WVOFF = 1.1883284e-08
+PVOFF = -9.6472405e-15
+NFACTOR = 1.247891
+LNFACTOR = -1.4165296e-07
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.03118654*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-4.3945878e-09*du0factorn_hp'
+WU0 = '-7.3769602e-10*du0factorn_hp'
+PU0 = '1.2865212e-15*du0factorn_hp'
+UA = 3.6660917e-27
+LUA = -6.37996e-34
+WUA = -2.2386272e-34
+PUA = 2.1442019e-40
+UB = 1e-19
+UC = -3.1451264e-27
+LUC = 1.7288353e-33
+WUC = 3.291833e-34
+PUC = -2.5730423e-40
+EU = 2.9
+VSAT = '108145.24*dvsatfactorn_hp'
+LVSAT = '-0.024092157*dvsatfactorn_hp'
+WVSAT = '-0.0014498529*dvsatfactorn_hp'
+PVSAT = '4.2884039e-09*dvsatfactorn_hp'
+A0 = 1.7986315
+LA0 = 5.9561165e-07
+WA0 = 8.6991173e-08
+PA0 = -2.5730423e-13
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5182587
+LUTE = -4.9634304e-08
+WUTE = 7.8877434e-09
+PUTE = 2.1442019e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.518 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.25303625+dvth0n518_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '5.4630255e-08+dlvth0n518_hp'
+WVTH0 = '-9.4607844e-09+dwvth0n518_hp'
+PVTH0 = '8.657897e-16+dpvth0n518_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14115967*dk2factorn_hp'
+LK2 = '-7.0826479e-09*dk2factorn_hp'
+WK2 = '-2.0373494e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11613396
+LVOFF = -2.430279e-08
+WVOFF = 6.6976194e-09
+PVOFF = -1.7283442e-15
+NFACTOR = 1.247891
+LNFACTOR = -1.4165296e-07
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.023930798*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '5.2650527e-09*du0factorn_hp'
+WU0 = '5.5382593e-10*du0factorn_hp'
+PU0 = '-4.3289485e-16*du0factorn_hp'
+UA = 3.3385821e-27
+LUA = 1.5394093e-33
+WUA = -1.6556601e-34
+PUA = -1.7315794e-40
+UB = 1e-19
+UC = -1.6439833e-27
+LUC = -4.0959891e-35
+WUC = 6.1979836e-35
+PUC = 5.7719314e-41
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2.287346
+LA0 = -8.4991775e-07
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.446538
+LUTE = -1.0239973e-08
+WUTE = -4.878535e-09
+PUTE = 1.4429828e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.618 NMOS
+LMIN = '1.00000000e-06+dlminn_hp'
+LMAX = '3.00000000e-06+dlmaxn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.25718806+dvth0n618_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.6064144e-08+dlvth0n618_hp'
+WVTH0 = '-9.8552056e-09+dwvth0n618_hp'
+PVTH0 = '3.5795702e-15+dpvth0n618_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.1583673*dk2factorn_hp'
+LK2 = '4.2495887e-08*dk2factorn_hp'
+WK2 = '-4.0262425e-10*dk2factorn_hp'
+PK2 = '-4.7099608e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.073115758
+LVOFF = -1.6172065e-08
+WVOFF = 2.6108905e-09
+PVOFF = -2.5007631e-15
+NFACTOR = 1.247891
+LNFACTOR = -1.4165296e-07
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.038208517*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.4279317e-08*du0factorn_hp'
+WU0 = '-8.0255738e-10*du0factorn_hp'
+PU0 = '2.3738203e-15*du0factorn_hp'
+UA = 3.9740572e-27
+LUA = -9.8023847e-33
+WUA = -2.2593614e-34
+PUA = 9.0431248e-40
+UB = 1e-19
+UC = -1.831564e-27
+LUC = 5.6661183e-34
+WUC = 7.98e-35
+PUC = 1.6896156e-56
+EU = 2.9
+VSAT = '173752.14*dvsatfactorn_hp'
+LVSAT = '-0.21814555*dvsatfactorn_hp'
+WVSAT = '-0.0070064533*dvsatfactorn_hp'
+PVSAT = '2.0723828e-08*dvsatfactorn_hp'
+A0 = 2.287346
+LA0 = -8.4991775e-07
+AGS = 0.452109
+LAGS = 1.4165296e-07
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.3407368
+LPCLM = 1.7528987e-07
+PDIBLC1 = 0
+PDIBLC2 = 0.0029224525
+LPDIBLC2 = 3.1871915e-09
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26991224
+LPVAG = -2.9318621e-08
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 4.005711e-09
+LALPHA0 = -2.9747121e-15
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.010447891
+LAIGC = -1.4165296e-10
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7049384
+LUTE = 3.399671e-07
+WUTE = 1.9669503e-08
+PUTE = -1.8839843e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.019 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '1.00000000e-05+dwminn0_hp'
+WMAX = '1.00000000e-04+wmaxoffsetn_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26788727+dvth0n019_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.1038171e-08+dlvth0n019_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.084018111
+LVOFF = -1.8808125e-11
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.035556364*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.0519085e-08*du0factorn_hp'
+UA = 3.7112729e-27
+LUA = -2.1038171e-33
+UB = 1e-19
+UC = -2.2112729e-27
+LUC = 2.1038171e-33
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+WVTH0 = '0.0+dwvth0n019_hp'
+PVTH0 = '0.0+dpvth0n019_hp'
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.119 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '3.00000000e-06+dwminn1_hp'
+WMAX = '1.00000000e-05+dwmaxn1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.26589897+dvth0n119_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.0001209e-08+dlvth0n119_hp'
+WVTH0 = '1.9739905e-08+dwvth0n119_hp'
+PVTH0 = '1.029496e-14+dpvth0n119_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.135*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.078708468
+LVOFF = -2.1381218e-09
+WVOFF = -5.2714141e-08
+PVOFF = 2.1040546e-14
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.035854024*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.1399508e-08*du0factorn_hp'
+WU0 = '-2.9551626e-09*du0factorn_hp'
+PU0 = '8.7408391e-15*du0factorn_hp'
+UA = 3.7996881e-27
+LUA = -2.98424e-33
+WUA = -8.7778641e-34
+PUA = 8.7408391e-39
+UB = 1e-19
+UC = -2.2112729e-27
+LUC = 2.1038171e-33
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.6911585
+LUTE = -8.8042295e-08
+WUTE = -8.7778641e-08
+PUTE = 8.7408391e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.219 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '1.00000000e-06+dwminn2_hp'
+WMAX = '3.00000000e-06+dwmaxn2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.27092513+dvth0n219_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '2.2513694e-08+dlvth0n219_hp'
+WVTH0 = '5.0182715e-09+dwvth0n219_hp'
+PVTH0 = '2.9358906e-15+dpvth0n219_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.12936476*dk2factorn_hp'
+LK2 = '-9.7876433e-09*dk2factorn_hp'
+WK2 = '-1.6505607e-08*dk2factorn_hp'
+PK2 = '2.8668007e-14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.083811759
+LVOFF = -5.5713177e-09
+WVOFF = -3.7766602e-08
+PVOFF = 3.1096377e-14
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.036402318*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.1645191e-08*du0factorn_hp'
+WU0 = '-4.5611173e-09*du0factorn_hp'
+PU0 = '9.4604423e-15*du0factorn_hp'
+UA = 3.5e-27
+UB = 1e-19
+UC = -2.3095639e-27
+LUC = 3.0825814e-33
+WUC = 2.8789441e-34
+PUC = -2.8668007e-39
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.7774796
+LUTE = 3.0825814e-07
+WUTE = 1.6505607e-07
+PUTE = -2.8668007e-13
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.319 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '5.00000000e-07+dwminn3_hp'
+WMAX = '1.00000000e-06+dwmaxn3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.28318117+dvth0n319_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '4.3867073e-08+dlvth0n319_hp'
+WVTH0 = '-6.3798453e-09+dwvth0n319_hp'
+PVTH0 = '-1.6922752e-14+dpvth0n319_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14986182*dk2factorn_hp'
+LK2 = '4.841314e-08*dk2factorn_hp'
+WK2 = '2.5566561e-09*dk2factorn_hp'
+PK2 = '-2.5458721e-14*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.11594168
+LVOFF = 1.1726934e-08
+WVOFF = -7.8857787e-09
+PVOFF = 1.5009003e-14
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.031813713*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.7248233e-09*du0factorn_hp'
+WU0 = '-2.9371434e-10*du0factorn_hp'
+PU0 = '-3.9036706e-15*du0factorn_hp'
+UA = 3.3533817e-27
+LUA = 1.4599984e-33
+WUA = 1.3635499e-34
+PUA = -1.3577985e-39
+UB = 1e-19
+UC = -2e-27
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.686747
+WUTE = 8.0674699e-08
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.419 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '2.40000000e-07+dwminn4_hp'
+WMAX = '5.00000000e-07+dwmaxn4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29237121+dvth0n419_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '3.7470129e-08+dlvth0n419_hp'
+WVTH0 = '-1.0349945e-08+dwvth0n419_hp'
+PVTH0 = '-1.4159272e-14+dpvth0n419_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.13619547*dk2factorn_hp'
+LK2 = '-1.7890728e-08*dk2factorn_hp'
+WK2 = '-3.3472055e-09*dk2factorn_hp'
+PK2 = '3.1845496e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.15520043
+LVOFF = 4.956697e-08
+WVOFF = 9.0740034e-09
+PVOFF = -1.337893e-15
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.031834606*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-6.3114512e-09*du0factorn_hp'
+WU0 = '-3.0274016e-10*du0factorn_hp'
+UA = 4.4181728e-27
+LUA = -2.8625165e-33
+WUA = -3.2363476e-34
+PUA = 5.0952793e-40
+UB = 1e-19
+UC = -2.3612495e-27
+LUC = -5.897314e-34
+WUC = 1.5605978e-34
+PUC = 2.5476397e-40
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5848845
+LUTE = 1.4743285e-07
+WUTE = 3.6670094e-08
+PUTE = -6.3690991e-14
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.519 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '1.50000000e-07+dwminn5_hp'
+WMAX = '2.40000000e-07+dwmaxn5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.29387256+dvth0n519_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '-6.6156176e-08+dlvth0n519_hp'
+WVTH0 = '-1.0617184e-08+dwvth0n519_hp'
+PVTH0 = '4.2862105e-15+dpvth0n519_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.14355422*dk2factorn_hp'
+WK2 = '-2.0373494e-09*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.13855729
+LVOFF = 4.2021388e-08
+WVOFF = 6.1115239e-09
+PVOFF = 5.2206043e-18
+NFACTOR = 1.2
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.030286984*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.3535401e-08*du0factorn_hp'
+WU0 = '-2.7263519e-11*du0factorn_hp'
+PU0 = '1.2858631e-15*du0factorn_hp'
+UA = 4.1846791e-27
+LUA = -9.6319336e-34
+WUA = -2.8207289e-34
+PUA = 1.7144842e-40
+UB = 1e-19
+UC = -2.2679835e-27
+LUC = 1.8047202e-33
+WUC = 1.3945843e-34
+PUC = -1.7144842e-40
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.3788727
+LUTE = -2.1038171e-07
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.MODEL NENHHP.619 NMOS
+LMIN = '3.00000000e-06+dlminn_hp'
+LMAX = '1.00000000e-05+lmaxoffsetn_hp'
+WMIN = '1.20000000e-07+wminoffsetn_hp'
+WMAX = '1.50000000e-07+dwmaxn6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.43e-09+dtoxn_hp'
+TOXP = '2.17e-09+dtoxn_hp'
+TOXM = 2.43e-09
+EPSROX = 3.9
+WINT = '3.59200000e-08+dwintn_hp'
+LINT = '2.10900000e-08+dlintn_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '2.75000000e-08+ddlcn_hp'
+DWC = '2.59200000e-08+ddwcn_hp'
+XPART = 0
+TOXREF = 2.43e-09
+DLCIG = 7.3824042e-09
+VTH0 = '0.22332363+dvth0n619_hp+(mcm_NENHHP_vth0*mcmScale)'
+LVTH0 = '1.2622902e-07+dlvth0n619_hp'
+WVTH0 = '-3.9150355e-09+dwvth0n619_hp'
+PVTH0 = '-1.3990384e-14+dpvth0n619_hp'
+K1 = '0.652*dk1factorn_hp'
+K2 = '-0.11412654*dk2factorn_hp'
+LK2 = '-8.8360317e-08*dk2factorn_hp'
+WK2 = '-4.8329787e-09*dk2factorn_hp'
+PK2 = '8.3942302e-15*dk2factorn_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.5e-08
+NGATE = 9e+21
+NDEP = 6.5e+17
+NSD = 1e+20
+PHIN = 5.960465e-09
+CDSC = 0
+CDSCB = -0.005
+CDSCD = 0
+CIT = 0
+VOFF = -0.058406899
+LVOFF = -5.9678222e-08
+WVOFF = -1.502763e-09
+PVOFF = 9.6666835e-15
+NFACTOR = 1.9966256
+LNFACTOR = -2.3562751e-06
+WNFACTOR = -7.5679432e-08
+PNFACTOR = 2.2384614e-13
+ETA0 = 0
+ETAB = -0.0731796
+U0 = '(0.03*du0factorn_hp)*(((1+mcm_NENHHP_u0*mcmScale)-1)+1)'
+UA = 7.7380366e-28
+LUA = -3.3661073e-34
+WUA = 4.1960284e-35
+PUA = 1.1192307e-40
+UB = 1e-19
+UC = -1.2416872e-27
+LUC = -1.1781376e-33
+WUC = 4.1960284e-35
+PUC = 1.1192307e-40
+EU = 2.9
+VSAT = '100000*dvsatfactorn_hp'
+A0 = 2
+AGS = 0.5
+A1 = 0
+A2 = 0.99
+B0 = 0
+B1 = 0
+KETA = 0.03
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 0.004
+PDIBLCB = 0.1
+DROUT = 0.56
+PVAG = 0.26
+DELTA = 0.01
+PSCBE1 = 2.882151e+09
+PSCBE2 = 0.00025
+FPROUT = 0
+PDITS = 0
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 144.8038
+RSW = 72.4019
+RDW = 72.4019
+PRWG = 0
+PRWB = 0.3
+WR = 1
+ALPHA0 = 1.1535274e-08
+LALPHA0 = -2.5245805e-14
+ALPHA1 = 3.309e-09
+BETA0 = 7
+AGIDL = 1.689e-07
+BGIDL = 2.879e+09
+CGIDL = 3.697
+EGIDL = -0.1135
+AIGBACC = 0.43
+BIGBACC = 0.054
+CIGBACC = 0.075
+NIGBACC = 0.5
+AIGBINV = 0.023
+BIGBINV = 0.008
+CIGBINV = 0.006
+EIGBINV = 1.1
+NIGBINV = 3
+AIGC = 0.0104
+BIGC = 0.001803274
+CIGC = 0.079999995
+AIGSD = 0.0086236294
+BIGSD = 0.00066508585
+CIGSD = 0.01875
+NIGC = 1
+POXEDGE = 1.105647
+PIGCD = 2.1
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1.01
+CGSO = '50.74e-12*dcgsofactorn_hp+dcgson_hp'
+CGDO = '50.74e-12*dcgdofactorn_hp+dcgdon_hp'
+CGBO = 0
+CGDL = '47.7e-12*dcgdlfactorn_hp'
+CGSL = '47.7e-12*dcgslfactorn_hp'
+CLC = 0
+CLE = 0.6
+CF = '135.61e-12*dcffactorn_hp'
+CKAPPAS = 0.9
+CKAPPAD = 0.9
+VFBCV = -0.8940079
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = 0
+KT1 = -0.1997
+KT1L = -1.4584643e-11
+KT2 = -0.03
+UTE = -1.5188727
+LUTE = -2.1038171e-07
+WUTE = 1.33e-08
+PUTE = 2.4851914e-28
+UA1 = 0
+UB1 = 0
+UC1 = 0
+PRT = 0
+AT = 50000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 1.5e-5
+JSWS = 3e-11
+JSWGS = 1e-07
+NJS = 1.54
+IJTHSFWD = 0.1
+JSD = 1.5e-5
+JSWD = 3e-11
+JSWGD = 1e-07
+NJD = 1.54
+IJTHDFWD = 0.1
+PBS = 729.7e-3
+CJS = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJS = 434.3e-3
+CJSWS = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWS = 193.6e-3
+PBSWGS = 1.170
+CJSWGS = '336.8e-12*dcjfactorn_hp'
+MJSWGS = 643.9e-3
+PBD = 729.7e-3
+CJD = '1.27e-3*dcjfactorn_hp+dcjn_hp'
+MJD = 434.3e-3
+PBSWD = 1.0
+CJSWD = '(43.24e-12-25e-9*1.27e-3)*dcjfactorn_hp'
+MJSWD = 193.6e-3
+PBSWGD = 1.170
+CJSWGD = '336.8e-12*dcjfactorn_hp'
+MJSWGD = 643.9e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjn_hp'
+XGW = 0
+XGL = 0
+RSHG = 8
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxln_hp'
+XW = '0.0+dxwn_hp'
+EM = 4.1e+07
+EF = 0.9
+NOIA = 8.25e+41
+NOIB = 1e+25
+NOIC = 8.75
+NTNOI = 1
+PBSWS = 1.0
+saref   = 2.43e-006       sbref   = 2.43e-006       wlod    = 0               kvth0   = 2.24e-009     
+lkvth0  = -2.67e-8        wkvth0  = -2.46e-10       pkvth0  = 0               llodvth = 3.33e-1             
+wlodvth = 3.33e-1         stk2    = 4e-10           lodk2   = 1               lodeta0 = 1             
+ku0     = -2.13e-9        lku0    = 1.26e-7         wku0    = 1.12e-7         pku0    = 0             
+llodku0 = 2.0e-1          wlodku0 = 2.0e-1          kvsat   = 0               steta0  = -4e-10             
+tku0    = 0             
+web     = 1.68e2          wec     = 1.88e3          kvth0we = 1.33e-2         k2we    = 0
+ku0we   = -9.35e-3        scref   = 1e-6            
+wpemod  = 1
.ENDS NENHHP_S


.SUBCKT PENHHP_S D G S B l=0 wpf=0 as=0 ad=0 ps=0 pd=0 nrs=0 nrd=0 simM=1 sa=0 sb=0 sc=0 sca=0 scb=0 scc=0 mcm_PENHHP_vth0=0 mcm_PENHHP_u0=0
** Pelgrom Scaling parameter **
.param mcmScale='1/sqrt(l*wpf)*1/sqrt(simM)'

.flat M0
M0 D G S B PENHHP l=l w=wpf as=as ad=ad ps=ps pd=pd nrs=nrs nrd=nrd
+ m=simM sa=sa sb=sb sc=sc sca=sca scb=scb scc=scc

.MODEL PENHHP.001 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p001_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.2243306
+NFACTOR = 0.9446555
+ETA0 = 0.3723176
+ETAB = -0.14
+U0 = '(0.0079*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1.8e-19
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 2.1
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.09
+DWG = 0
+DWB = 0
+PCLM = 1.4
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p001_hp'
+WVTH0 = '0.0+dwvth0p001_hp'
+PVTH0 = '0.0+dpvth0p001_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.101 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38424489+dvth0p101_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '4.2321575e-08+dwvth0p101_hp'
+K1 = '0.65424489*dk1factorp_hp'
+WK1 = '-4.2321575e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.20692654
+WVOFF = -1.7351846e-07
+NFACTOR = 0.73241089
+WNFACTOR = 2.1160787e-06
+ETA0 = 0.3723176
+ETAB = -0.13575511
+WETAB = -4.2321575e-08
+U0 = '(0.0077302043*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '1.692863e-09*du0factorp_hp'
+UA = 1.8848978e-19
+WUA = -8.4643149e-26
+UB = 1e-19
+UC = -1.1273468e-19
+WUC = 1.2696472e-25
+EU = 2
+VSAT = '161510.22*dvsatfactorp_hp'
+WVSAT = '0.084643149*dvsatfactorp_hp'
+A0 = 2.1848978
+WA0 = -8.4643149e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.094244892
+WKETA = -4.2321575e-08
+DWG = 0
+DWB = 0
+PCLM = 1.3151022
+WPCLM = 8.4643149e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p101_hp'
+PVTH0 = '0.0+dpvth0p101_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.201 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.36270635+dvth0p201_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '-2.1669425e-08+dwvth0p201_hp'
+K1 = '0.64*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.25317452
+WVOFF = -3.6115708e-08
+NFACTOR = 1.3960312
+WNFACTOR = 1.4446283e-07
+ETA0 = 0.36745517
+WETA0 = 1.4446283e-08
+ETAB = -0.15972486
+WETAB = 2.8892566e-08
+U0 = '(0.0084458729*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-4.3338849e-10*du0factorp_hp'
+UA = 1.2596298e-19
+WUA = 1.0112398e-25
+UB = 1e-19
+UC = -6.5137569e-20
+WUC = -1.4446283e-26
+EU = 2
+VSAT = '194862.43*dvsatfactorp_hp'
+WVSAT = '-0.014446283*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p201_hp'
+PVTH0 = '0.0+dpvth0p201_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.301 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.40879518+dvth0p301_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '2.3128916e-08+dwvth0p301_hp'
+K1 = '0.64951807*dk1factorp_hp'
+WK1 = '-9.2515663e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.35981253
+WVOFF = 6.7536434e-08
+NFACTOR = 1.9253784
+WNFACTOR = -3.7006265e-07
+ETA0 = 0.47749832
+WETA0 = -9.2515663e-08
+ETAB = -0.12048193
+WETAB = -9.2515663e-09
+U0 = '(0.0082855422*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-2.7754699e-10*du0factorp_hp'
+UA = 1.4433735e-19
+WUA = 8.3264096e-26
+UB = 1e-19
+UC = -6.0963855e-20
+WUC = -1.8503133e-26
+EU = 2
+VSAT = '180000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.8855422
+WPCLM = -2.7754699e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p301_hp'
+PVTH0 = '0.0+dpvth0p301_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.401 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.33401575+dvth0p401_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '-1.2316535e-08+dwvth0p401_hp'
+K1 = '0.64732283*dk1factorp_hp'
+WK1 = '-8.2110236e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.20607076
+WVOFF = -5.3371654e-09
+NFACTOR = 1.1446555
+ETA0 = 0.26499477
+WETA0 = 8.2110236e-09
+ETAB = -0.13133858
+WETAB = -4.1055118e-09
+U0 = '(0.0072669291*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '2.0527559e-10*du0factorp_hp'
+UA = 3.719685e-19
+WUA = -2.4633071e-26
+UB = 1e-19
+UC = -1.1732283e-19
+WUC = 8.2110236e-27
+EU = 2
+VSAT = '180000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.3866142
+WPCLM = -4.1055118e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p401_hp'
+PVTH0 = '0.0+dpvth0p401_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.501 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.47253012+dvth0p501_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '1.8156627e-08+dwvth0p501_hp'
+K1 = '0.6760241*dk1factorp_hp'
+WK1 = '-1.4525301e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.31286072
+WVOFF = 1.8156627e-08
+NFACTOR = 0.48441454
+WNFACTOR = 1.4525301e-07
+ETA0 = 0.50038989
+WETA0 = -4.3575904e-08
+ETAB = -0.19951807
+WETAB = 1.0893976e-08
+U0 = '(0.0083650602*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-3.6313253e-11*du0factorp_hp'
+UA = 2.9301205e-19
+WUA = -7.2626506e-27
+UB = 1e-19
+UC = -9.6506024e-20
+WUC = 3.6313253e-27
+EU = 2
+VSAT = '196506.02*dvsatfactorp_hp'
+WVSAT = '-0.0036313253*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 0.86987952
+WPCLM = 7.2626506e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p501_hp'
+PVTH0 = '0.0+dpvth0p501_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.601 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.34+dvth0p601_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.4804*dk1factorp_hp'
+WK1 = '1.22752e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1579306
+WVOFF = -3.0688e-09
+NFACTOR = 1.9926555
+WNFACTOR = -6.1376e-08
+ETA0 = 0.0927176
+WETA0 = 1.22752e-08
+ETAB = -0.0752
+WETAB = -6.1376e-09
+U0 = '(0.00586*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.0688e-10*du0factorp_hp'
+UA = 8.672e-19
+WUA = -8.59264e-26
+UB = 1e-19
+UC = -2.52e-20
+WUC = -6.1376e-27
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = -0.392
+WPCLM = 2.45504e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0071246
+WAIGC = 6.44448e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p601_hp'
+WVTH0 = '0.0+dwvth0p601_hp'
+PVTH0 = '0.0+dpvth0p601_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.701 PMOS
+LMIN = '9.19000000e-08+lminoffsetp_hp'
+LMAX = '9.44500000e-08+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.34+dvth0p701_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.59*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1853306
+NFACTOR = 1.4446555
+ETA0 = 0.2023176
+ETAB = -0.13
+U0 = '(0.0086*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1e-19
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.8
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 5.2e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p701_hp'
+WVTH0 = '0.0+dwvth0p701_hp'
+PVTH0 = '0.0+dpvth0p701_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.002 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p002_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.0292534
+LVOFF = -1.3300481e-08
+NFACTOR = -1.8729445
+LNFACTOR = 1.4778312e-07
+ETA0 = 0.0905576
+LETA0 = 1.4778312e-08
+ETAB = -0.23392
+LETAB = 4.926104e-09
+U0 = '(0.0060216*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '9.852208e-11*du0factorp_hp'
+UA = 1.8e-19
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '357840*dvsatfactorp_hp'
+LVSAT = '-0.009852208*dvsatfactorp_hp'
+A0 = 1.1608
+LA0 = 4.926104e-08
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.00392
+LKETA = 4.926104e-09
+DWG = 0
+DWB = 0
+PCLM = 3.2784
+LPCLM = -9.852208e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p002_hp'
+WVTH0 = '0.0+dwvth0p002_hp'
+PVTH0 = '0.0+dpvth0p002_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.102 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.34437687+dvth0p102_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.091078e-09+dlvth0p102_hp'
+WVTH0 = '-3.5516265e-07+dwvth0p102_hp'
+PVTH0 = '2.0848048e-14+dpvth0p102_hp'
+K1 = '0.61437687*dk1factorp_hp'
+LK1 = '2.091078e-09*dk1factorp_hp'
+WK1 = '3.5516265e-07*dk1factorp_hp'
+PK1 = '-2.0848048e-14*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.076933426
+LVOFF = -6.818139e-09
+WVOFF = 1.0586827e-06
+PVOFF = -6.4628948e-14
+NFACTOR = -0.091787763
+LNFACTOR = 4.322922e-08
+WNFACTOR = -1.7758133e-05
+PNFACTOR = 1.0424024e-12
+ETA0 = 0.0905576
+LETA0 = 1.4778312e-08
+ETAB = -0.26954313
+LETAB = 7.017182e-09
+WETAB = 3.5516265e-07
+PETAB = -2.0848048e-14
+U0 = '(0.0074465254*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.487896e-11*du0factorp_hp'
+WU0 = '-1.4206506e-08*du0factorp_hp'
+PU0 = '8.3392191e-16*du0factorp_hp'
+UA = 1.0875373e-19
+LUA = 4.182156e-27
+WUA = 7.1032531e-25
+PUA = -4.1696095e-32
+UB = 1e-19
+UC = 6.8694042e-21
+LUC = -6.273234e-27
+WUC = -1.065488e-24
+PUC = 6.2544143e-32
+EU = 2
+VSAT = '429086.27*dvsatfactorp_hp'
+LVSAT = '-0.014034364*dvsatfactorp_hp'
+WVSAT = '-0.71032531*dvsatfactorp_hp'
+PVSAT = '4.1696095e-08*dvsatfactorp_hp'
+A0 = 0.84701757
+LA0 = 7.017182e-08
+WA0 = 3.1284108e-06
+PA0 = -2.0848048e-13
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.039543135
+LKETA = 7.017182e-09
+WKETA = 3.5516265e-07
+PKETA = -2.0848048e-14
+DWG = 0
+DWB = 0
+PCLM = 3.9908627
+LPCLM = -1.4034364e-07
+WPCLM = -7.1032531e-06
+PPCLM = 4.1696095e-13
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.202 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.52512828+dvth0p202_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '8.5190303e-09+dlvth0p202_hp'
+WVTH0 = '1.8184981e-07+dwvth0p202_hp'
+PVTH0 = '-1.0674584e-14+dpvth0p202_hp'
+K1 = '0.73392*dk1factorp_hp'
+LK1 = '-4.926104e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.086055685
+LVOFF = -1.7792624e-08
+WVOFF = 5.74442e-07
+PVOFF = -3.2023752e-14
+NFACTOR = -5.6608893
+LNFACTOR = 3.7013548e-07
+WNFACTOR = -1.2123321e-06
+PNFACTOR = 7.1163893e-14
+ETA0 = 0.13136312
+LETA0 = 1.2383028e-08
+WETA0 = -1.2123321e-07
+PETA0 = 7.1163893e-15
+ETAB = -0.068388954
+LETAB = -4.7905684e-09
+WETAB = -2.4246642e-07
+PETAB = 1.4232779e-14
+U0 = '(0.0014406343*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.6742477e-10*du0factorp_hp'
+WU0 = '3.6369962e-09*du0factorp_hp'
+PU0 = '-2.1349168e-16*du0factorp_hp'
+UA = 2.6813503e-19
+LUA = -7.4569238e-27
+WUA = 2.3680347e-25
+PUA = -7.1163893e-33
+UB = 1e-19
+UC = -3.9256552e-19
+LUC = 1.7173596e-26
+WUC = 1.2123321e-25
+PUC = -7.1163893e-33
+EU = 2
+VSAT = '149194.48*dvsatfactorp_hp'
+LVSAT = '0.0023952842*dvsatfactorp_hp'
+WVSAT = '0.12123321*dvsatfactorp_hp'
+PVSAT = '-7.1163893e-09*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.302 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.13835084+dvth0p302_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.4184805e-08+dlvth0p302_hp'
+WVTH0 = '-1.9409786e-07+dwvth0p302_hp'
+PVTH0 = '1.1393544e-14+dpvth0p302_hp'
+K1 = '0.83283181*dk1factorp_hp'
+LK1 = '-9.6148054e-09*dk1factorp_hp'
+WK1 = '-9.6142277e-08*dk1factorp_hp'
+PK1 = '4.5574178e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 1.170744
+LVOFF = -8.027769e-08
+WVOFF = -4.7987504e-07
+PVOFF = 2.8711732e-14
+NFACTOR = -10.103171
+LNFACTOR = 6.3089742e-07
+WNFACTOR = 3.1055658e-06
+PNFACTOR = -1.8229671e-13
+ETA0 = -0.52393782
+LETA0 = 5.2525326e-08
+WETA0 = 5.1571931e-07
+PETA0 = -3.1901924e-14
+ETAB = -0.39771566
+LETAB = 1.4540909e-08
+WETAB = 7.7639144e-08
+PETAB = -4.5574178e-15
+U0 = '(0.0036800675*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.4155715e-10*du0factorp_hp'
+WU0 = '1.4602672e-09*du0factorp_hp'
+PU0 = '-9.1148355e-17*du0factorp_hp'
+UA = 6.9427855e-19
+LUA = -2.8844416e-26
+WUA = -1.7740803e-25
+PUA = 1.3672253e-32
+UB = 1e-19
+UC = -4.2759133e-19
+LUC = 1.9229611e-26
+WUC = 1.5527829e-25
+PUC = -9.1148355e-33
+EU = 2
+VSAT = '363313.73*dvsatfactorp_hp'
+LVSAT = '-0.0096148054*dvsatfactorp_hp'
+WVSAT = '-0.08689071*dvsatfactorp_hp'
+PVSAT = '4.5574178e-09*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.8855422
+WPCLM = -2.7754699e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.402 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.84724787+dvth0p402_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '2.6919025e-08+dlvth0p402_hp'
+WVTH0 = '1.4191933e-07+dwvth0p402_hp'
+PVTH0 = '-8.0896713e-15+dpvth0p402_hp'
+K1 = '0.5659748*dk1factorp_hp'
+LK1 = '4.2667043e-09*dk1factorp_hp'
+WK1 = '3.0347943e-08*dk1factorp_hp'
+PK1 = '-2.0224178e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.088261211
+LVOFF = -1.5437712e-08
+WVOFF = 3.3221802e-08
+PVOFF = -2.0224178e-15
+NFACTOR = -3.5513445
+LNFACTOR = 2.463052e-07
+ETA0 = 0.79079886
+LETA0 = -2.7578425e-08
+WETA0 = -1.0746588e-07
+PETA0 = 6.0672534e-15
+ETAB = -0.30660661
+LETAB = 9.1928083e-09
+WETAB = 3.4453455e-08
+PETAB = -2.0224178e-15
+U0 = '(0.0079546898*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.6073045e-11*du0factorp_hp'
+WU0 = '-5.6590375e-10*du0factorp_hp'
+PU0 = '4.0448356e-17*du0factorp_hp'
+UA = 2.0927244e-19
+LUA = 8.5334085e-27
+WUA = 5.2484863e-26
+PUA = -4.0448356e-33
+UB = 1e-19
+UC = 4.5373228e-20
+LUC = -8.5334085e-27
+WUC = -6.890691e-26
+PUC = 4.0448356e-33
+EU = 2
+VSAT = '180000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.3866142
+WPCLM = -4.1055118e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.502 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '0.56794506+dvth0p502_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.4572923e-08+dlvth0p502_hp'
+WVTH0 = '-1.6942311e-07+dwvth0p502_hp'
+PVTH0 = '9.8385574e-15+dpvth0p502_hp'
+K1 = '0.61491952*dk1factorp_hp'
+LK1 = '3.2049351e-09*dk1factorp_hp'
+WK1 = '1.9580106e-08*dk1factorp_hp'
+PK1 = '-1.7888286e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.77683759
+LVOFF = -5.7154677e-08
+WVOFF = -1.18265e-07
+PVOFF = 7.1553144e-15
+NFACTOR = 1.9893977
+LNFACTOR = -7.8936365e-08
+WNFACTOR = -1.2189633e-06
+PNFACTOR = 7.1553144e-14
+ETA0 = -1.3599051
+LETA0 = 9.757247e-08
+WETA0 = 3.6568898e-07
+PETA0 = -2.1465943e-14
+ETAB = 0.26555566
+LETAB = -2.4393117e-08
+WETAB = -9.1422246e-08
+PETAB = 5.3664858e-15
+U0 = '(0.0039972145*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.2909351e-10*du0factorp_hp'
+WU0 = '3.0474082e-10*du0factorp_hp'
+PU0 = '-1.7888286e-17*du0factorp_hp'
+UA = 1.7080289e-19
+LUA = 6.4098703e-27
+WUA = 6.0948164e-26
+PUA = -3.5776572e-33
+UB = 1e-19
+UC = -1.2932145e-19
+LUC = 1.7211689e-27
+WUC = -3.0474082e-26
+PUC = 1.7888286e-33
+EU = 2
+VSAT = '196506.02*dvsatfactorp_hp'
+WVSAT = '-0.0036313253*dvsatfactorp_hp'
+A0 = 1.1248771
+LA0 = 4.0655196e-08
+WA0 = 1.7052704e-07
+PA0 = -8.944143e-15
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 3.9703711
+LPCLM = -1.6262078e-07
+WPCLM = -6.0948164e-07
+PPCLM = 3.5776572e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.19899508
+LKT1 = -1.6262078e-09
+WKT1 = -6.8210814e-09
+PKT1 = 3.5776572e-16
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.602 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-1.2998624+dvth0p602_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '5.0344783e-08+dlvth0p602_hp'
+WVTH0 = '8.6466509e-08+dwvth0p602_hp'
+PVTH0 = '-4.5351684e-15+dpvth0p602_hp'
+K1 = '1.5097632*dk1factorp_hp'
+LK1 = '-5.39901e-08*dk1factorp_hp'
+WK1 = '-1.0301348e-07*dk1factorp_hp'
+PK1 = '6.0468912e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.9055338
+LVOFF = 3.9211788e-08
+WVOFF = 1.1221988e-07
+PVOFF = -6.0468912e-15
+NFACTOR = -10.667761
+LNFACTOR = 6.6403882e-07
+WNFACTOR = 5.1506739e-07
+PNFACTOR = -3.0234456e-14
+ETA0 = 2.0612808
+LETA0 = -1.0325114e-07
+WETA0 = -1.0301348e-07
+PETA0 = 6.0468912e-15
+ETAB = -0.7777216
+LETAB = 3.6847258e-08
+WETAB = 5.1506739e-08
+PETAB = -3.0234456e-15
+U0 = '(0.016604448*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-5.635463e-10*du0factorp_hp'
+WU0 = '-1.4224502e-09*du0factorp_hp'
+PU0 = '9.0703368e-17*du0factorp_hp'
+UA = 2.9259264e-18
+LUA = -1.079802e-25
+WUA = -3.1650376e-25
+PUA = 1.2093782e-32
+UB = 1e-19
+UC = -7.277216e-19
+LUC = 3.6847258e-26
+WUC = 5.1506739e-26
+PUC = -3.0234456e-33
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 4.473408
+LA0 = -1.3497525e-07
+WA0 = -2.882217e-07
+PA0 = 1.5117228e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.937216
+LPCLM = -1.2216738e-07
+WPCLM = -3.3093939e-07
+PPCLM = 3.0234456e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0071246
+WAIGC = 6.44448e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = 0.21405376
+LKT1 = -2.329062e-08
+WKT1 = -6.3408773e-08
+PKT1 = 3.3257902e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.702 PMOS
+LMIN = '9.44500000e-08+dlminp_hp'
+LMAX = '1.00700000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.52784+dvth0p702_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '9.852208e-09+dlvth0p702_hp'
+K1 = '0.59*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.0964294
+LVOFF = -1.4778312e-08
+NFACTOR = -6.0689445
+LNFACTOR = 3.9408832e-07
+ETA0 = 1.1415176
+LETA0 = -4.926104e-08
+ETAB = -0.31784
+LETAB = 9.852208e-09
+U0 = '(0.003904*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.463052e-10*du0factorp_hp'
+UA = 1e-19
+UB = 1e-19
+UC = -2.6784e-19
+LUC = 9.852208e-27
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = -1.0176
+LPCLM = 1.4778312e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.086032e-07
+LALPHA0 = 8.4236378e-15
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.352096
+LKT1 = 6.4039352e-09
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p702_hp'
+PVTH0 = '0.0+dpvth0p702_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.003 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p003_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1973306
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.0077*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1.8e-19
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 2
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.49e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p003_hp'
+WVTH0 = '0.0+dwvth0p003_hp'
+PVTH0 = '0.0+dpvth0p003_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.103 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p103_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.19308571
+WVOFF = -4.2321575e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.0077*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1.8e-19
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 2.0424489
+WA0 = -4.2321575e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.49e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p103_hp'
+WVTH0 = '0.0+dwvth0p103_hp'
+PVTH0 = '0.0+dpvth0p103_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.203 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p203_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.21705546
+WVOFF = 2.8892566e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.0077*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1.4110055e-19
+WUA = 1.1557027e-25
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.49e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p203_hp'
+WVTH0 = '0.0+dwvth0p203_hp'
+PVTH0 = '0.0+dpvth0p203_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.303 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p303_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.19684867
+WVOFF = 9.2515663e-09
+NFACTOR = 0.6446555
+ETA0 = 0.37087182
+WETA0 = -2.7754699e-08
+ETAB = -0.15
+U0 = '(0.0077951807*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-9.2515663e-11*du0factorp_hp'
+UA = 2.0289157e-19
+WUA = 5.5509398e-26
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '199518.07*dvsatfactorp_hp'
+WVSAT = '-0.0092515663*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.8855422
+WPCLM = -2.7754699e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.49e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p303_hp'
+WVTH0 = '0.0+dwvth0p303_hp'
+PVTH0 = '0.0+dpvth0p303_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.403 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38866142+dvth0p403_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '4.1055118e-09+dwvth0p403_hp'
+K1 = '0.63866142*dk1factorp_hp'
+WK1 = '-4.1055118e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.17473217
+WVOFF = -1.2316535e-09
+NFACTOR = 0.6446555
+ETA0 = 0.32097902
+WETA0 = -4.1055118e-09
+ETAB = -0.15
+U0 = '(0.0073401575*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '1.2316535e-10*du0factorp_hp'
+UA = 3.5464567e-19
+WUA = -1.6422047e-26
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '180000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.3866142
+WPCLM = -4.1055118e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.49e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007595
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p403_hp'
+PVTH0 = '0.0+dpvth0p403_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.503 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.62523751+dvth0p503_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '1.5466894e-08+dlvth0p503_hp'
+WVTH0 = '5.6152252e-08+dwvth0p503_hp'
+PVTH0 = '-3.4027166e-15+dpvth0p503_hp'
+K1 = '0.77491422*dk1factorp_hp'
+LK1 = '-6.1867537e-09*dk1factorp_hp'
+WK1 = '-3.4081128e-08*dk1factorp_hp'
+PK1 = '1.3610858e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.46032714
+LVOFF = 1.5466894e-08
+WVOFF = 6.159924e-08
+PVOFF = -3.4027166e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0068460386*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '6.1867537e-11*du0factorp_hp'
+WU0 = '2.3187152e-10*du0factorp_hp'
+PU0 = '-1.3610858e-17*du0factorp_hp'
+UA = 8.0698136e-19
+LUA = -3.0933806e-26
+WUA = -1.159359e-25
+PUA = 6.8054373e-33
+UB = 1e-19
+UC = -3.1079254e-19
+LUC = 1.2373522e-26
+WUC = 4.637436e-26
+PUC = -2.7221749e-33
+EU = 2
+VSAT = '196506.02*dvsatfactorp_hp'
+WVSAT = '-0.0036313253*dvsatfactorp_hp'
+A0 = 2.3444522
+LA0 = -3.0933862e-08
+WA0 = -9.7779483e-08
+PA0 = 6.8054496e-15
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = -0.90792608
+LPCLM = 1.2373526e-07
+WPCLM = 4.6374374e-07
+PPCLM = -2.7221757e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.6965962e-07
+LALPHA0 = -1.965039e-14
+WALPHA0 = -7.3647116e-14
+PALPHA0 = 4.3230857e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0075423014
+LAIGC = 3.0934049e-12
+WAIGC = 1.1593681e-11
+PAIGC = -6.8054909e-19
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2477779
+LKT1 = 1.2373432e-09
+WKT1 = 3.9111372e-09
+PKT1 = -2.7221551e-16
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.603 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '0.43258853+dvth0p603_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.1350087e-08+dlvth0p603_hp'
+WVTH0 = '-8.8769915e-08+dwvth0p603_hp'
+PVTH0 = '5.7512097e-15+dpvth0p603_hp'
+K1 = '0.2400848*dk1factorp_hp'
+LK1 = '2.0540022e-08*dk1factorp_hp'
+WK1 = '3.9190502e-08*dk1factorp_hp'
+PK1 = '-2.3004825e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.63725793
+LVOFF = -5.1350087e-08
+WVOFF = -8.8769915e-08
+PVOFF = 5.7512097e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.010503152*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0540022e-10*du0factorp_hp'
+WU0 = '-2.6915302e-10*du0factorp_hp'
+PU0 = '2.3004825e-17*du0factorp_hp'
+UA = -6.6317811e-19
+LUA = 1.0270024e-25
+WUA = 8.5475949e-26
+PUA = -1.1502426e-32
+UB = 1e-19
+UC = 5.9983125e-19
+LUC = -4.1080094e-26
+WUC = -7.8381099e-26
+PUC = 4.6009705e-33
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 0.42441871
+LA0 = 1.0270042e-07
+WA0 = 1.652651e-07
+PA0 = -1.1502447e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 6.8543146
+LPCLM = -4.1080107e-07
+WPCLM = -5.9968323e-07
+PPCLM = 4.6009719e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -1.0765019e-06
+LALPHA0 = 6.5239294e-14
+WALPHA0 = 1.2447702e-13
+PALPHA0 = -7.3068009e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0072995592
+LAIGC = -1.0270104e-11
+WAIGC = 4.4849371e-11
+PAIGC = 1.1502517e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.11273738
+LKT1 = -4.1079795e-09
+WKT1 = -1.4589413e-08
+PKT1 = 4.6009371e-16
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.703 PMOS
+LMIN = '1.00700000e-07+dlminp_hp'
+LMAX = '1.03900000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.36+dvth0p703_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.59*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1553306
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0081*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1e-19
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.5
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.49e-08
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.243
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p703_hp'
+WVTH0 = '0.0+dwvth0p703_hp'
+PVTH0 = '0.0+dpvth0p703_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.004 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p004_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.016551379
+LVOFF = -1.1190234e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.010411688*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.6785351e-10*du0factorp_hp'
+UA = 8.961039e-20
+LUA = 5.5951169e-27
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 1.0961039
+LA0 = 5.5951169e-08
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.19116883
+LKETA = 1.6785351e-08
+DWG = 0
+DWB = 0
+PCLM = 2.5038961
+LPCLM = -5.5951169e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -2.5219548e-07
+LALPHA0 = 1.777121e-14
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076401948
+LAIGC = -2.7975584e-12
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p004_hp'
+WVTH0 = '0.0+dwvth0p004_hp'
+PVTH0 = '0.0+dpvth0p004_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.104 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p104_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.012306487
+LVOFF = -1.1190234e-08
+WVOFF = -4.2321575e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.011179077*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.1535484e-10*du0factorp_hp'
+WU0 = '-7.6508613e-09*du0factorp_hp'
+PU0 = '4.7358831e-16*du0factorp_hp'
+UA = 5.1240975e-20
+LUA = 7.9701836e-27
+WUA = 3.8254306e-25
+PUA = -2.3679416e-32
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 0.75485867
+LA0 = 7.9701836e-08
+WA0 = 3.4022149e-06
+PA0 = -2.3679416e-13
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.19116883
+LKETA = 1.6785351e-08
+DWG = 0
+DWB = 0
+PCLM = 2.5038961
+LPCLM = -5.5951169e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -2.5219548e-07
+LALPHA0 = 1.777121e-14
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076401948
+LAIGC = -2.7975584e-12
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p104_hp'
+WVTH0 = '0.0+dwvth0p104_hp'
+PVTH0 = '0.0+dpvth0p104_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.204 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.42395133+dvth0p204_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '2.7205871e-09+dlvth0p204_hp'
+WVTH0 = '1.3057939e-07+dwvth0p204_hp'
+PVTH0 = '-8.0828643e-15+dpvth0p204_hp'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.036276242
+LVOFF = -1.1190234e-08
+WVOFF = 2.8892566e-08
+PVOFF = -2.2434455e-29
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.0090434094*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-8.315704e-11*du0factorp_hp'
+WU0 = '-1.3057939e-09*du0factorp_hp'
+PU0 = '8.0828643e-17*du0factorp_hp'
+UA = 1.4110055e-19
+WUA = 1.1557027e-25
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.19116883
+LKETA = 1.6785351e-08
+DWG = 0
+DWB = 0
+PCLM = 2.9434094
+LPCLM = -8.315704e-08
+WPCLM = -1.3057939e-06
+PPCLM = 8.0828643e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -2.5219548e-07
+LALPHA0 = 1.777121e-14
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076401948
+LAIGC = -2.7975584e-12
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.304 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.30925553+dvth0p304_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-4.3790825e-09+dlvth0p304_hp'
+WVTH0 = '1.909508e-08+dwvth0p304_hp'
+PVTH0 = '-1.1819854e-15+dpvth0p304_hp'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.10315825
+LVOFF = -1.8570428e-08
+WVOFF = -1.0663776e-07
+PVOFF = 7.1735491e-15
+NFACTOR = 0.6446555
+ETA0 = 0.37087182
+WETA0 = -2.7754699e-08
+ETAB = -0.15
+U0 = '(0.0051532154*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6353765e-10*du0factorp_hp'
+WU0 = '2.4754746e-09*du0factorp_hp'
+PU0 = '-1.589586e-16*du0factorp_hp'
+UA = 2.5573084e-19
+LUA = -3.2707509e-27
+WUA = 4.1496259e-27
+PUA = 3.1791699e-33
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '146678.8*dvsatfactorp_hp'
+LVSAT = '0.0032707509*dvsatfactorp_hp'
+WVSAT = '0.042108205*dvsatfactorp_hp'
+PVSAT = '-3.1791699e-09*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.29075139
+LKETA = 2.2949511e-08
+WKETA = 9.6794251e-08
+PKETA = -5.9915641e-15
+DWG = 0
+DWB = 0
+PCLM = 0.30036317
+LPCLM = 9.812258e-08
+WPCLM = 1.263247e-06
+PPCLM = -9.5375148e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -3.5762686e-07
+LALPHA0 = 2.4297412e-14
+WALPHA0 = 1.024793e-13
+PALPHA0 = -6.3434686e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076832115
+LAIGC = -5.4602948e-12
+WAIGC = -4.1812274e-11
+PAIGC = 2.5881797e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.404 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.25975495+dvth0p404_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-7.9793103e-09+dlvth0p404_hp'
+WVTH0 = '-4.3681967e-09+dwvth0p404_hp'
+PVTH0 = '5.2452256e-16+dpvth0p404_hp'
+K1 = '0.75609674*dk1factorp_hp'
+LK1 = '-7.2692463e-09*dk1factorp_hp'
+WK1 = '-5.9769854e-08*dk1factorp_hp'
+PK1 = '3.4456228e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.22771435
+LVOFF = 3.2795964e-09
+WVOFF = 5.0195853e-08
+PVOFF = -3.1833626e-15
+NFACTOR = 0.6446555
+ETA0 = 0.32097902
+WETA0 = -4.1055118e-09
+ETAB = -0.15
+U0 = '(0.012520074*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.2063681e-10*du0factorp_hp'
+WU0 = '-1.0164162e-09*du0factorp_hp'
+PU0 = '7.0540099e-17*du0factorp_hp'
+UA = 2.5104741e-19
+LUA = 6.4127321e-27
+WUA = 6.3695691e-27
+PUA = -1.4108011e-33
+UB = 1e-19
+UC = -2.5658043e-19
+LUC = 9.6923285e-27
+WUC = 7.4219123e-26
+PUC = -4.5941637e-33
+EU = 2
+VSAT = '283598.26*dvsatfactorp_hp'
+LVSAT = '-0.0064127321*dvsatfactorp_hp'
+WVSAT = '-0.022791616*dvsatfactorp_hp'
+PVSAT = '1.4108011e-09*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.0040757206
+LKETA = 4.6997129e-09
+WKETA = -4.2953801e-08
+PKETA = 2.6588403e-15
+DWG = 0
+DWB = 0
+PCLM = 2.1458571
+LPCLM = -4.6997139e-08
+WPCLM = 3.8848286e-07
+PPCLM = -2.6588401e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -4.5483568e-08
+LALPHA0 = 4.9757429e-15
+WALPHA0 = -4.5476621e-14
+PALPHA0 = 2.8150028e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0075558549
+LAIGC = 2.4230821e-12
+WAIGC = 1.8554781e-11
+PAIGC = -1.1485409e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.504 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38565079+dvth0p504_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '6.3647549e-10+dlvth0p504_hp'
+WVTH0 = '2.3328887e-08+dwvth0p504_hp'
+PVTH0 = '-1.3709503e-15+dpvth0p504_hp'
+K1 = '0.41553401*dk1factorp_hp'
+LK1 = '1.6058881e-08*dk1factorp_hp'
+WK1 = '1.5153947e-08*dk1factorp_hp'
+PK1 = '-1.6865653e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.018846496
+LVOFF = -1.4193955e-08
+WVOFF = -4.0475326e-09
+PVOFF = 6.6081863e-16
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0068460369*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '6.1867642e-11*du0factorp_hp'
+WU0 = '2.3187189e-10*du0factorp_hp'
+PU0 = '-1.3610881e-17*du0factorp_hp'
+UA = 8.069813e-19
+LUA = -3.0933802e-26
+WUA = -1.1593589e-25
+PUA = 6.8054365e-33
+UB = 1e-19
+UC = 1.6838132e-19
+LUC = -1.728734e-26
+WUC = -1.9272461e-26
+PUC = 1.3413633e-33
+EU = 2
+VSAT = '196506.02*dvsatfactorp_hp'
+WVSAT = '-0.0036313253*dvsatfactorp_hp'
+A0 = 2.3444508
+LA0 = -3.0933775e-08
+WA0 = -9.7779173e-08
+PA0 = 6.8054304e-15
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.63876076
+LKETA = 4.4491291e-08
+WKETA = 9.8470224e-08
+PKETA = -6.0953069e-15
+DWG = 0
+DWB = 0
+PCLM = 6.2796826
+LPCLM = -3.2117772e-07
+WPCLM = -5.2095875e-07
+PPCLM = 3.3731327e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -3.9131636e-07
+LALPHA0 = 2.7454024e-14
+WALPHA0 = 3.0606594e-14
+PALPHA0 = -2.1302189e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076620955
+LAIGC = -4.3218469e-12
+WAIGC = -4.8181532e-12
+PAIGC = 3.3534347e-19
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.24777811
+LKT1 = 1.2373565e-09
+WKT1 = 3.9111844e-09
+PKT1 = -2.7221844e-16
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.604 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '0.43258918+dvth0p604_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.1350127e-08+dlvth0p604_hp'
+WVTH0 = '-8.8769989e-08+dwvth0p604_hp'
+PVTH0 = '5.7512142e-15+dpvth0p604_hp'
+K1 = '1.0499751*dk1factorp_hp'
+LK1 = '-2.959219e-08*dk1factorp_hp'
+WK1 = '-7.1764489e-08*dk1factorp_hp'
+PK1 = '4.5676315e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.63725858
+LVOFF = -5.1350127e-08
+WVOFF = -8.8769989e-08
+PVOFF = 5.7512142e-15
+NFACTOR = 0.6446555
+ETA0 = 1.1122085
+LETA0 = -5.0132247e-08
+WETA0 = -1.1095505e-07
+PETA0 = 6.8681179e-15
+ETAB = -0.15
+U0 = '(-0.025941933*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.0505506e-09*du0factorp_hp'
+WU0 = '4.7238238e-09*du0factorp_hp'
+PU0 = '-2.8606044e-16*du0factorp_hp'
+UA = -6.6317793e-19
+LUA = 1.0270022e-25
+WUA = 8.5475928e-26
+PUA = -1.1502425e-32
+UB = 1e-19
+UC = -2.1005974e-19
+LUC = 9.0521578e-27
+WUC = 3.2573963e-26
+PUC = -2.2671479e-33
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 0.42442339
+LA0 = 1.0270013e-07
+WA0 = 1.6526458e-07
+PA0 = -1.1502415e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 6.8543108
+LPCLM = -4.1080083e-07
+WPCLM = -5.9968281e-07
+PPCLM = 4.6009693e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 2.0968584e-07
+LALPHA0 = -1.437573e-14
+WALPHA0 = -5.1730708e-14
+PALPHA0 = 3.6004573e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.011349012
+LAIGC = -2.6093122e-10
+WAIGC = -5.0992568e-10
+PAIGC = 3.5490827e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.63916576
+LKT1 = 2.8477937e-08
+WKT1 = 5.7531293e-08
+PKT1 = -4.004178e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.704 PMOS
+LMIN = '1.03900000e-07+dlminp_hp'
+LMAX = '1.11600000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.36+dvth0p704_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.40922078*dk1factorp_hp'
+LK1 = '1.1190234e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1553306
+NFACTOR = 0.6446555
+ETA0 = 0.12153838
+LETA0 = 1.1190234e-08
+ETAB = -0.15
+U0 = '(0.016235065*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-5.0356052e-10*du0factorp_hp'
+UA = 1e-19
+UB = 1e-19
+UC = 8.0779221e-20
+LUC = -1.1190234e-26
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.5
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -2.5219548e-07
+LALPHA0 = 1.777121e-14
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0067961039
+LAIGC = 5.5951169e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.12549351
+LKT1 = -7.2736519e-09
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p704_hp'
+WVTH0 = '0.0+dwvth0p704_hp'
+PVTH0 = '0.0+dpvth0p704_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.005 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p005_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1773306
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.008*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1.7e-19
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 1.7
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p005_hp'
+WVTH0 = '0.0+dwvth0p005_hp'
+PVTH0 = '0.0+dpvth0p005_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.105 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38+dvth0p105_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.17308571
+WVOFF = -4.2321575e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.0080848978*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-8.4643149e-10*du0factorp_hp'
+UA = 1.6575511e-19
+WUA = 4.2321575e-26
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 1.7
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p105_hp'
+WVTH0 = '0.0+dwvth0p105_hp'
+PVTH0 = '0.0+dpvth0p105_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.205 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38486243+dvth0p205_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '1.4446283e-08+dwvth0p205_hp'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.19705546
+WVOFF = 2.8892566e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3423176
+ETAB = -0.15
+U0 = '(0.0078486243*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-1.4446283e-10*du0factorp_hp'
+UA = 1.4110055e-19
+WUA = 1.1557027e-25
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '190000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 1.7486243
+WPCLM = -1.4446283e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p205_hp'
+PVTH0 = '0.0+dpvth0p205_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.305 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.46616048+dvth0p305_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '6.541502e-09+dlvth0p305_hp'
+WVTH0 = '9.3467989e-08+dwvth0p305_hp'
+PVTH0 = '-6.3583399e-15+dpvth0p305_hp'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.21065186
+LVOFF = 3.2707552e-09
+WVOFF = 4.2108266e-08
+PVOFF = -3.1791741e-15
+NFACTOR = 0.6446555
+ETA0 = 0.37087182
+WETA0 = -2.7754699e-08
+ETAB = -0.15
+U0 = '(0.0051532163*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.6353759e-10*du0factorp_hp'
+WU0 = '2.4754738e-09*du0factorp_hp'
+PU0 = '-1.5895854e-16*du0factorp_hp'
+UA = 2.557309e-19
+LUA = -3.2707552e-27
+WUA = 4.1495652e-27
+PUA = 3.1791741e-33
+UB = 1e-19
+UC = -1e-19
+EU = 2
+VSAT = '146678.74*dvsatfactorp_hp'
+LVSAT = '0.0032707552*dvsatfactorp_hp'
+WVSAT = '0.042108266*dvsatfactorp_hp'
+PVSAT = '-3.1791741e-09*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.17996368
+LKETA = -9.8122581e-09
+WKETA = -1.263247e-07
+PKETA = 9.5375149e-15
+DWG = 0
+DWB = 0
+PCLM = 0.30036328
+LPCLM = 9.8122572e-08
+WPCLM = 1.2632469e-06
+PPCLM = -9.537514e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 1.4073488e-07
+LALPHA0 = -1.0388565e-14
+WALPHA0 = -1.3374417e-13
+PALPHA0 = 1.0097685e-20
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0075438595
+LAIGC = 4.2386073e-12
+WAIGC = 5.456856e-11
+PAIGC = -4.1199263e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.405 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.1901263+dvth0p405_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.2825465e-08+dlvth0p405_hp'
+WVTH0 = '-3.7372215e-08+dwvth0p405_hp'
+PVTH0 = '2.8216022e-15+dpvth0p405_hp'
+K1 = '0.65165354*dk1factorp_hp'
+WK1 = '-1.026378e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.088456631
+LVOFF = -6.4127406e-09
+WVOFF = -1.5812273e-08
+PVOFF = 1.4108029e-15
+NFACTOR = 0.6446555
+ETA0 = 0.32097902
+WETA0 = -4.1055118e-09
+ETAB = -0.15
+U0 = '(0.012520072*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-3.206367e-10*du0factorp_hp'
+WU0 = '-1.0164158e-09*du0factorp_hp'
+PU0 = '7.0540073e-17*du0factorp_hp'
+UA = 2.5104729e-19
+LUA = 6.4127406e-27
+WUA = 6.3695961e-27
+PUA = -1.4108029e-33
+UB = 1e-19
+UC = -1.1732283e-19
+WUC = 8.2110236e-27
+EU = 2
+VSAT = '283598.38*dvsatfactorp_hp'
+LVSAT = '-0.0064127406*dvsatfactorp_hp'
+WVSAT = '-0.022791643*dvsatfactorp_hp'
+PVSAT = '1.4108029e-09*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.20481069
+LKETA = 1.9238207e-08
+WKETA = 5.6058351e-08
+PKETA = -4.2324055e-15
+DWG = 0
+DWB = 0
+PCLM = 4.2347208
+LPCLM = -1.9238205e-07
+WPCLM = -6.0163858e-07
+PPCLM = 4.2324051e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = -2.6663856e-07
+LALPHA0 = 2.0368131e-14
+WALPHA0 = 5.9350844e-14
+PALPHA0 = -4.4809887e-21
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077100707
+LAIGC = -8.3103403e-12
+WAIGC = -2.4215561e-11
+PAIGC = 1.8282749e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.505 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.37650602+dvth0p505_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '3.6313253e-09+dwvth0p505_hp'
+K1 = '0.64626506*dk1factorp_hp'
+WK1 = '-9.0783133e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.18508964
+WVOFF = 5.446988e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0077349398*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.6313253e-11*du0factorp_hp'
+UA = 3.6253012e-19
+WUA = -1.8156627e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '196506.02*dvsatfactorp_hp'
+WVSAT = '-0.0036313253*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.00048192771
+WKETA = 1.0893976e-08
+DWG = 0
+DWB = 0
+PCLM = 1.6650602
+WPCLM = -3.6313253e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p505_hp'
+PVTH0 = '0.0+dpvth0p505_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.605 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.3052+dvth0p605_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '-6.1376e-09+dwvth0p605_hp'
+K1 = '0.6248*dk1factorp_hp'
+WK1 = '-6.1376e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1005306
+WVOFF = -6.1376e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3919176
+WETA0 = -1.22752e-08
+ETAB = -0.15
+U0 = '(0.00352*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '6.1376e-10*du0factorp_hp'
+UA = 8.124e-19
+WUA = -7.97888e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 0.952
+WPCLM = 6.1376e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p605_hp'
+PVTH0 = '0.0+dpvth0p605_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.705 PMOS
+LMIN = '1.11600000e-07+dlminp_hp'
+LMAX = '1.17500000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.36+dvth0p705_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.57*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1553306
+NFACTOR = 0.6446555
+ETA0 = 0.2823176
+ETAB = -0.15
+U0 = '(0.009*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 1e-19
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '170000*dvsatfactorp_hp'
+A0 = 1.9
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.5
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p705_hp'
+WVTH0 = '0.0+dwvth0p705_hp'
+PVTH0 = '0.0+dpvth0p705_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.006 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32097403+dvth0p006_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-4.456461e-09+dlvth0p006_hp'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.00025267792
+LVOFF = -1.3369383e-08
+NFACTOR = 0.6446555
+ETA0 = 0.5784215
+LETA0 = -1.7825844e-08
+ETAB = -0.15
+U0 = '(0.0068194805*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.9129221e-11*du0factorp_hp'
+UA = 7.6025974e-19
+LUA = -4.456461e-26
+UB = 1e-19
+UC = -2.7707792e-19
+LUC = 1.3369383e-26
+EU = 2
+VSAT = '249025.97*dvsatfactorp_hp'
+LVSAT = '-0.004456461*dvsatfactorp_hp'
+A0 = 0.12922078
+LA0 = 1.3369383e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 2.2902597
+LPCLM = -4.456461e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0084853896
+LAIGC = -6.6846916e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0056293912
+LAIGSD = 3.1195227e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 5.9025974e-19
+LUC1 = -4.456461e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p006_hp'
+PVTH0 = '0.0+dpvth0p006_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.106 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.34602992+dvth0p106_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.5647414e-09+dlvth0p106_hp'
+WVTH0 = '2.4980722e-07+dwvth0p106_hp'
+PVTH0 = '-1.8860445e-14+dpvth0p106_hp'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.021063675
+LVOFF = -1.1477663e-08
+WVOFF = 2.0748564e-07
+PVOFF = -1.8860445e-14
+NFACTOR = 0.6446555
+ETA0 = 0.5784215
+LETA0 = -1.7825844e-08
+ETAB = -0.15
+U0 = '(0.0064032606*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.2696361e-10*du0factorp_hp'
+WU0 = '4.1497128e-09*du0factorp_hp'
+PU0 = '-3.772089e-16*du0factorp_hp'
+UA = 8.3118252e-19
+LUA = -5.0239769e-26
+WUA = -7.0710007e-25
+PUA = 5.6581334e-32
+UB = 1e-19
+UC = -3.0213381e-19
+LUC = 1.5261103e-26
+WUC = 2.4980722e-25
+PUC = -1.8860445e-32
+EU = 2
+VSAT = '249025.97*dvsatfactorp_hp'
+LVSAT = '-0.004456461*dvsatfactorp_hp'
+A0 = -0.12133811
+LA0 = 1.5261103e-07
+WA0 = 2.4980722e-06
+PA0 = -1.8860445e-13
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 2.2902597
+LPCLM = -4.456461e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0084853896
+LAIGC = -6.6846916e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.005454
+LAIGSD = 4.4437265e-11
+WAIGSD = 1.7486505e-09
+PAIGSD = -1.3202311e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 8.4081863e-19
+LUC1 = -6.3481807e-26
+WUC1 = -2.4980721e-24
+PUC1 = 1.8860445e-31
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.206 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.23810951+dvth0p206_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.1079846e-08+dlvth0p206_hp'
+WVTH0 = '-7.082431e-08+dwvth0p206_hp'
+PVTH0 = '6.4379298e-15+dpvth0p206_hp'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.10506067
+LVOFF = -2.2809768e-08
+WVOFF = -1.672298e-07
+PVOFF = 1.4807239e-14
+NFACTOR = 0.6446555
+ETA0 = 0.63582344
+LETA0 = -2.2159691e-08
+WETA0 = -1.7054119e-07
+PETA0 = 1.287586e-14
+ETAB = -0.15
+U0 = '(0.0078486243*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-1.4446283e-10*du0factorp_hp'
+UA = 6.1168432e-19
+LUA = -3.5529074e-26
+WUA = -5.4970922e-26
+PUA = 1.287586e-32
+UB = 1e-19
+UC = -2.1805195e-19
+LUC = 8.9129221e-27
+EU = 2
+VSAT = '263376.46*dvsatfactorp_hp'
+LVSAT = '-0.0055399228*dvsatfactorp_hp'
+WVSAT = '-0.042635297*dvsatfactorp_hp'
+PVSAT = '3.2189649e-09*dvsatfactorp_hp'
+A0 = 1.0064903
+LA0 = 6.7459986e-08
+WA0 = -8.5270593e-07
+PA0 = 6.4379298e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 2.0518743
+LPCLM = -2.2895375e-08
+WPCLM = 7.082431e-07
+PPCLM = -6.4379298e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0084853896
+LAIGC = -6.6846916e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.17259805
+LKT1 = -4.3338471e-09
+WKT1 = -1.7054119e-07
+PKT1 = 1.287586e-14
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.306 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.3204921+dvth0p306_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-4.456461e-09+dlvth0p306_hp'
+WVTH0 = '9.2515663e-09+dwvth0p306_hp'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.083840849
+LVOFF = -6.3034762e-09
+WVOFF = 1.6382481e-08
+PVOFF = -1.2368773e-15
+NFACTOR = 0.6446555
+ETA0 = 0.60128646
+LETA0 = -1.7396306e-08
+WETA0 = -1.3697124e-07
+PETA0 = 8.2458489e-15
+ETAB = -0.15
+U0 = '(0.0073192771*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.7006265e-10*du0factorp_hp'
+UA = 6.1990221e-19
+LUA = -3.0765689e-26
+WUA = -6.2958711e-26
+PUA = 8.2458489e-33
+UB = 1e-19
+UC = -2.1805195e-19
+LUC = 8.9129221e-27
+EU = 2
+VSAT = '247603.66*dvsatfactorp_hp'
+LVSAT = '-0.0043490764*dvsatfactorp_hp'
+WVSAT = '-0.027304136*dvsatfactorp_hp'
+PVSAT = '2.0614622e-09*dvsatfactorp_hp'
+A0 = -0.43259271
+LA0 = 1.7611075e-07
+WA0 = 5.4608271e-07
+PA0 = -4.1229245e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.10618135
+LKETA = -4.2416918e-09
+WKETA = -5.4608271e-08
+PKETA = 4.1229245e-15
+DWG = 0
+DWB = 0
+PCLM = 3.9041465
+LPCLM = -1.7396306e-07
+WPCLM = -1.0921654e-06
+PPCLM = 8.2458489e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0084853896
+LAIGC = -6.6846916e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.46041465
+LKT1 = 1.7396306e-08
+WKT1 = 1.0921654e-07
+PKT1 = -8.2458489e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+PVTH0 = '0.0+dpvth0p306_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.406 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.30097403+dvth0p406_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-4.456461e-09+dlvth0p406_hp'
+K1 = '0.65165354*dk1factorp_hp'
+WK1 = '-1.026378e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.014441757
+LVOFF = -1.2000864e-08
+WVOFF = -1.6512688e-08
+PVOFF = 1.4636843e-15
+NFACTOR = 0.6446555
+ETA0 = 0.32097902
+WETA0 = -4.1055118e-09
+ETAB = -0.15
+U0 = '(0.0082732283*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-8.2110236e-11*du0factorp_hp'
+UA = 6.6643675e-19
+LUA = -2.4949164e-26
+WUA = -8.5016085e-26
+PUA = 5.488816e-33
+UB = 1e-19
+UC = -3.376245e-19
+LUC = 1.6632776e-26
+WUC = 5.667739e-26
+PUC = -3.6592107e-33
+EU = 2
+VSAT = '121974.13*dvsatfactorp_hp'
+LVSAT = '0.0057898903*dvsatfactorp_hp'
+WVSAT = '0.032244263*dvsatfactorp_hp'
+PVSAT = '-2.744408e-09*dvsatfactorp_hp'
+A0 = 1.2307291
+LA0 = 5.0529952e-08
+WA0 = -2.4233183e-07
+PA0 = 1.8296053e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.060150833
+LKETA = 8.3163879e-09
+WKETA = 2.4233183e-08
+PKETA = -1.8296053e-15
+DWG = 0
+DWB = 0
+PCLM = 1.6866142
+WPCLM = -4.1055118e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0084853896
+LAIGC = -6.6846916e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0053399794
+LAIGSD = 5.3045817e-11
+WAIGSD = 3.3302937e-10
+PAIGSD = -2.5143717e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p406_hp'
+PVTH0 = '0.0+dpvth0p406_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.506 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.41490847+dvth0p506_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '2.8993843e-09+dlvth0p506_hp'
+WVTH0 = '2.5065577e-08+dwvth0p506_hp'
+PVTH0 = '-1.618286e-15+dpvth0p506_hp'
+K1 = '0.74369348*dk1factorp_hp'
+LK1 = '-7.3558453e-09*dk1factorp_hp'
+WK1 = '-3.0512565e-08*dk1factorp_hp'
+PK1 = '1.618286e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.094772784
+LVOFF = -6.8189223e-09
+WVOFF = 1.1601377e-09
+PVOFF = 3.2365719e-16
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0077349398*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.6313253e-11*du0factorp_hp'
+UA = 3.6253012e-19
+WUA = -1.8156627e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '431187.61*dvsatfactorp_hp'
+LVSAT = '-0.01771846*dvsatfactorp_hp'
+WVSAT = '-0.035782702*dvsatfactorp_hp'
+PVSAT = '2.427429e-09*dvsatfactorp_hp'
+A0 = -2.7936317
+LA0 = 3.5436919e-07
+WA0 = 6.4302754e-07
+PA0 = -4.8548579e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.19533876
+LKETA = -1.4711691e-08
+WKETA = -3.1974527e-08
+PKETA = 3.2365719e-15
+DWG = 0
+DWB = 0
+PCLM = 1.6650602
+WPCLM = -3.6313253e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0109211
+LAIGC = -2.5074305e-10
+WAIGC = -5.3585628e-10
+PAIGC = 4.0457149e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0042955421
+LAIGSD = 1.3190083e-10
+WAIGSD = 5.6280557e-10
+PAIGSD = -4.249182e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.52228524
+LKT1 = 2.2067536e-08
+WKT1 = 6.4302754e-08
+PKT1 = -4.8548579e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.606 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.05492987+dvth0p606_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.8895395e-08+dlvth0p606_hp'
+WVTH0 = '-2.4251491e-08+dwvth0p606_hp'
+PVTH0 = '1.3675988e-15+dpvth0p606_hp'
+K1 = '0.30133766*dk1factorp_hp'
+LK1 = '2.4421406e-08*dk1factorp_hp'
+WK1 = '3.0090182e-08*dk1factorp_hp'
+PK1 = '-2.7351975e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.049437717
+LVOFF = -3.8575127e-09
+WVOFF = -5.0507665e-09
+PVOFF = -8.2055926e-17
+NFACTOR = 0.6446555
+ETA0 = 0.3919176
+WETA0 = -1.22752e-08
+ETAB = -0.15
+U0 = '(-0.0044130909*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '5.9894836e-10*du0factorp_hp'
+WU0 = '1.7005935e-09*du0factorp_hp'
+PU0 = '-8.2055926e-17*du0factorp_hp'
+UA = 2.9278909e-18
+LUA = -1.5971956e-25
+WUA = -3.6961105e-25
+PUA = 2.188158e-32
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '-94436.364*dvsatfactorp_hp'
+LVSAT = '0.019964945*dvsatfactorp_hp'
+WVSAT = '0.036227782*dvsatfactorp_hp'
+PVSAT = '-2.7351975e-09*dvsatfactorp_hp'
+A0 = 7.1887273
+LA0 = -3.9929891e-07
+WA0 = -7.2455564e-07
+PA0 = 5.4703951e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.56692468
+LKETA = 4.8842813e-08
+WKETA = 7.2455564e-08
+PKETA = -5.4703951e-15
+DWG = 0
+DWB = 0
+PCLM = -1.6923636
+LPCLM = 1.9964945e-07
+WPCLM = 4.2365382e-07
+PPCLM = -2.7351975e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0096541039
+LAIGC = -1.5508484e-10
+WAIGC = -3.6227782e-10
+PAIGC = 2.7351975e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.008403612
+LAIGSD = -1.7825844e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -1.3751039
+LKT1 = 8.6455344e-08
+WKT1 = 1.8113891e-07
+PKT1 = -1.3675988e-14
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = -2.6443636e-18
+LUC1 = 1.9964945e-25
+WUC1 = 3.6227782e-25
+PUC1 = -2.7351975e-32
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.706 PMOS
+LMIN = '1.17500000e-07+dlminp_hp'
+LMAX = '1.32900000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.27146104+dvth0p706_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-6.6846916e-09+dlvth0p706_hp'
+K1 = '0.57*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.094533847
+LVOFF = -4.5901549e-09
+NFACTOR = 0.6446555
+ETA0 = 0.2823176
+ETAB = -0.15
+U0 = '(0.010770779*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.3369383e-10*du0factorp_hp'
+UA = -3.7220779e-19
+LUA = 3.5651688e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '229025.97*dvsatfactorp_hp'
+LVSAT = '-0.004456461*dvsatfactorp_hp'
+A0 = 0.71948052
+LA0 = 8.9129221e-08
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 2.0902597
+LPCLM = -4.456461e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0064194805
+LAIGC = 8.9129221e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.008403612
+LAIGSD = -1.7825844e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = 0.24220779
+LKT1 = -3.5651688e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 5.9025974e-19
+LUC1 = -4.456461e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p706_hp'
+PVTH0 = '0.0+dpvth0p706_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.007 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.37+dvth0p007_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1473306
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0078*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 2.7e-19
+UB = 1e-19
+UC = -1.3e-19
+EU = 2
+VSAT = '200000*dvsatfactorp_hp'
+A0 = 1.6
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 1.8
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.005972573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-19
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p007_hp'
+WVTH0 = '0.0+dwvth0p007_hp'
+PVTH0 = '0.0+dpvth0p007_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.107 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.37424489+dvth0p107_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '4.2321575e-08+dwvth0p107_hp'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1473306
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0078*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 2.7848978e-19
+WUA = -8.4643149e-26
+UB = 1e-19
+UC = -1.3424489e-19
+WUC = 4.2321575e-26
+EU = 2
+VSAT = '200000*dvsatfactorp_hp'
+A0 = 1.5575511
+WA0 = 4.2321575e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 1.8
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0059428588
+WAIGSD = 2.9625102e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.4244892e-19
+WUC1 = -4.2321574e-25
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p107_hp'
+PVTH0 = '0.0+dpvth0p107_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.207 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.36+dvth0p207_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.14587187
+WVOFF = -4.3338849e-09
+NFACTOR = 0.6446555
+ETA0 = 0.39204246
+WETA0 = -2.8892566e-08
+ETAB = -0.15
+U0 = '(0.0078486243*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-1.4446283e-10*du0factorp_hp'
+UA = 2.2082541e-19
+WUA = 8.6677699e-26
+UB = 1e-19
+UC = -1.2e-19
+EU = 2
+VSAT = '202431.22*dvsatfactorp_hp'
+WVSAT = '-0.0072231416*dvsatfactorp_hp'
+A0 = 1.7486243
+WA0 = -1.4446283e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.05
+DWG = 0
+DWB = 0
+PCLM = 1.8
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.22027514
+WKT1 = -2.8892566e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p207_hp'
+WVTH0 = '0.0+dwvth0p207_hp'
+PVTH0 = '0.0+dpvth0p207_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.307 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.36951807+dvth0p307_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '9.2515663e-09+dwvth0p307_hp'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.15318602
+WVOFF = 2.7754699e-09
+NFACTOR = 0.6446555
+ETA0 = 0.40990796
+WETA0 = -4.6257831e-08
+ETAB = -0.15
+U0 = '(0.0073192771*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.7006265e-10*du0factorp_hp'
+UA = 2.8144578e-19
+WUA = 2.7754699e-26
+UB = 1e-19
+UC = -1.2e-19
+EU = 2
+VSAT = '199759.04*dvsatfactorp_hp'
+WVSAT = '-0.0046257831*dvsatfactorp_hp'
+A0 = 1.5048193
+WA0 = 9.2515663e-08
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.059518072
+WKETA = -9.2515663e-09
+DWG = 0
+DWB = 0
+PCLM = 1.9903614
+WPCLM = -1.8503133e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.26903614
+WKT1 = 1.8503133e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p307_hp'
+PVTH0 = '0.0+dpvth0p307_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.407 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.35+dvth0p407_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.65165354*dk1factorp_hp'
+WK1 = '-1.026378e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.14646446
+WVOFF = -4.1055118e-10
+NFACTOR = 0.6446555
+ETA0 = 0.32097902
+WETA0 = -4.1055118e-09
+ETAB = -0.15
+U0 = '(0.0082732283*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '-8.2110236e-11*du0factorp_hp'
+UA = 3.919685e-19
+WUA = -2.4633071e-26
+UB = 1e-19
+UC = -1.5464567e-19
+WUC = 1.6422047e-26
+EU = 2
+VSAT = '185669.29*dvsatfactorp_hp'
+WVSAT = '0.0020527559*dvsatfactorp_hp'
+A0 = 1.7866142
+WA0 = -4.1055118e-08
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.031338583
+WKETA = 4.1055118e-09
+DWG = 0
+DWB = 0
+PCLM = 1.6866142
+WPCLM = -4.1055118e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0059235417
+WAIGSD = 5.6420817e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p407_hp'
+WVTH0 = '0.0+dwvth0p407_hp'
+PVTH0 = '0.0+dpvth0p407_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.507 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.38301205+dvth0p507_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '7.2626506e-09+dwvth0p507_hp'
+K1 = '0.66277108*dk1factorp_hp'
+WK1 = '-1.2709639e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.16978843
+WVOFF = 4.7207229e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0077349398*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.6313253e-11*du0factorp_hp'
+UA = 3.6253012e-19
+WUA = -1.8156627e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '236265.06*dvsatfactorp_hp'
+WVSAT = '-0.0090783133*dvsatfactorp_hp'
+A0 = 1.1048193
+WA0 = 1.0893976e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.033493976
+WKETA = 3.6313253e-09
+DWG = 0
+DWB = 0
+PCLM = 1.6650602
+WPCLM = -3.6313253e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0081626506
+WAIGC = -9.0783133e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0057465964
+WAIGSD = 9.5348798e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.27951807
+WKT1 = 1.0893976e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p507_hp'
+PVTH0 = '0.0+dpvth0p507_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.607 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.2628+dvth0p607_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '-9.2064e-09+dwvth0p607_hp'
+K1 = '0.57*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.0918746
+WVOFF = -5.953472e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3919176
+WETA0 = -1.22752e-08
+ETAB = -0.15
+U0 = '(0.002176*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '7.97888e-10*du0factorp_hp'
+UA = 1.1708e-18
+WUA = -1.288896e-25
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '125200*dvsatfactorp_hp'
+WVSAT = '0.0061376*dvsatfactorp_hp'
+A0 = 2.796
+WA0 = -1.22752e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.0296
+WKETA = 1.22752e-08
+DWG = 0
+DWB = 0
+PCLM = 0.504
+WPCLM = 1.22752e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007948
+WAIGC = -6.1376e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006442573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.424
+WKT1 = 3.0688e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = -4.48e-19
+WUC1 = 6.1376e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p607_hp'
+PVTH0 = '0.0+dpvth0p607_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.707 PMOS
+LMIN = '1.32900000e-07+dlminp_hp'
+LMAX = '1.38700000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.345+dvth0p707_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.57*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1450306
+NFACTOR = 0.6446555
+ETA0 = 0.2823176
+ETAB = -0.15
+U0 = '(0.0093*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 2e-20
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '180000*dvsatfactorp_hp'
+A0 = 1.7
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0074
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006442573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-19
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p707_hp'
+WVTH0 = '0.0+dwvth0p707_hp'
+PVTH0 = '0.0+dpvth0p707_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.008 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.29173045+dvth0p008_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-7.5686656e-09+dlvth0p008_hp'
+K1 = '0.67608985*dk1factorp_hp'
+LK1 = '-2.5228885e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.0951509
+LVOFF = -5.045777e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0075391015*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.5228885e-11*du0factorp_hp'
+UA = 4.5262895e-19
+LUA = -1.766022e-26
+UB = 1e-19
+UC = -1.0391015e-19
+LUC = -2.5228885e-27
+EU = 2
+VSAT = '239134.78*dvsatfactorp_hp'
+LVSAT = '-0.0037843328*dvsatfactorp_hp'
+A0 = 0.29550749
+LA0 = 1.2614443e-07
+AGS = -0.11391015
+LAGS = -2.5228885e-09
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.054359401
+LKETA = 1.0091554e-08
+DWG = 0
+DWB = 0
+PCLM = 2.321797
+LPCLM = -5.045777e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006155202
+LAIGSD = -1.766022e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = -1.608985e-19
+LUC1 = 2.5228885e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p008_hp'
+PVTH0 = '0.0+dpvth0p008_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.108 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.28490048+dvth0p108_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-8.6396045e-09+dlvth0p108_hp'
+WVTH0 = '-6.809478e-08+dwvth0p108_hp'
+PVTH0 = '1.0677261e-14+dpvth0p108_hp'
+K1 = '0.67608985*dk1factorp_hp'
+LK1 = '-2.5228885e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.0951509
+LVOFF = -5.045777e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0075391015*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '2.5228885e-11*du0factorp_hp'
+UA = 4.3896902e-19
+LUA = -1.5518342e-26
+WUA = 1.3618956e-25
+PUA = -2.1354523e-32
+UB = 1e-19
+UC = -9.7080182e-20
+LUC = -3.5938275e-27
+WUC = -6.809478e-26
+PUC = 1.0677261e-32
+EU = 2
+VSAT = '239134.78*dvsatfactorp_hp'
+LVSAT = '-0.0037843328*dvsatfactorp_hp'
+A0 = 0.36380717
+LA0 = 1.1543504e-07
+WA0 = -6.809478e-07
+PA0 = 1.0677261e-13
+AGS = -0.12498501
+LAGS = -1.4519496e-09
+WAGS = 1.1041635e-07
+PAGS = -1.0677261e-14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.054359401
+LKETA = 1.0091554e-08
+DWG = 0
+DWB = 0
+PCLM = 2.4325456
+LPCLM = -6.116716e-08
+WPCLM = -1.1041635e-06
+PPCLM = 1.0677261e-13
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006150487
+LAIGSD = -2.007765e-11
+WAIGSD = 4.7008185e-11
+PAIGSD = 2.4101782e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -0.98322458
+LUTE = 3.2128169e-09
+WUTE = 3.3124906e-07
+PUTE = -3.2031784e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = -2.2919818e-19
+LUC1 = 3.5938275e-26
+WUC1 = 6.8094779e-25
+PUC1 = -1.0677261e-31
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.208 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.3078203+dvth0p208_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.045777e-09+dlvth0p208_hp'
+K1 = '0.68877586*dk1factorp_hp'
+LK1 = '-3.7496257e-09*dk1factorp_hp'
+WK1 = '-3.7690136e-08*dk1factorp_hp'
+PK1 = '3.6446362e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.089886367
+LVOFF = -5.4137982e-09
+WVOFF = -1.5640926e-08
+PVOFF = 1.0933909e-15
+NFACTOR = 0.6446555
+ETA0 = 0.36667044
+LETA0 = 2.4534744e-09
+WETA0 = 4.6487706e-08
+PETA0 = -7.2892724e-15
+ETAB = -0.15
+U0 = '(0.0074608657*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.7496257e-11*du0factorp_hp'
+WU0 = '2.3243853e-10*du0factorp_hp'
+PU0 = '-3.6446362e-17*du0factorp_hp'
+UA = 5.3175013e-19
+LUA = -3.006642e-26
+WUA = -1.3946312e-25
+PUA = 2.1867817e-32
+UB = 1e-19
+UC = -1.2e-19
+EU = 2
+VSAT = '247909*dvsatfactorp_hp'
+LVSAT = '-0.0043977014*dvsatfactorp_hp'
+WVSAT = '-0.02606821*dvsatfactorp_hp'
+PVSAT = '1.8223181e-09*dvsatfactorp_hp'
+A0 = -0.19734701
+LA0 = 1.8817543e-07
+WA0 = 9.8624126e-07
+PA0 = -1.0933909e-13
+AGS = -0.062448279
+LAGS = -7.4992514e-09
+WAGS = -7.5380273e-08
+PAGS = 7.2892724e-15
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.054359401
+LKETA = 1.0091554e-08
+DWG = 0
+DWB = 0
+PCLM = 2.0608985
+LPCLM = -2.5228885e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0061663093
+LAIGSD = -1.1965303e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.24564716
+LKT1 = 2.4534744e-09
+WKT1 = 4.6487706e-08
+PKT1 = -7.2892724e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.83367242
+LUTE = -1.1248877e-08
+WUTE = -1.1307041e-07
+PUTE = 1.0933909e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p208_hp'
+PVTH0 = '0.0+dpvth0p208_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.308 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.29250586+dvth0p308_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-7.4470806e-09+dlvth0p308_hp'
+WVTH0 = '-1.4885632e-08+dwvth0p308_hp'
+PVTH0 = '2.334067e-15+dpvth0p308_hp'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.091450521
+LVOFF = -5.969823e-09
+WVOFF = -1.4120569e-08
+PVOFF = 1.6338469e-15
+NFACTOR = 0.6446555
+ETA0 = 0.33792512
+LETA0 = 6.9607406e-09
+WETA0 = 7.4428158e-08
+PETA0 = -1.1670335e-14
+ETAB = -0.15
+U0 = '(0.0083125774*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-9.6052141e-11*du0factorp_hp'
+WU0 = '-5.9542526e-10*du0factorp_hp'
+PU0 = '9.3362681e-17*du0factorp_hp'
+UA = 3.8454784e-19
+LUA = -9.9699691e-27
+WUA = 3.617501e-27
+PUA = 2.334067e-33
+UB = 1e-19
+UC = -1.2e-19
+EU = 2
+VSAT = '213432.63*dvsatfactorp_hp'
+LVSAT = '-0.0013222368*dvsatfactorp_hp'
+WVSAT = '0.0074428158*dvsatfactorp_hp'
+PVSAT = '-1.1670335e-09*dvsatfactorp_hp'
+A0 = 1.2187739
+LA0 = 2.7660585e-08
+WA0 = -3.9022829e-07
+PA0 = 4.6681341e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.044841329
+LKETA = 1.0091554e-08
+WKETA = -9.2515663e-09
+PKETA = -4.0489609e-31
+DWG = 0
+DWB = 0
+PCLM = 1.5062847
+LPCLM = 4.6810221e-08
+WPCLM = 5.3908461e-07
+PPCLM = -7.0022011e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0062840825
+LAIGSD = -2.3353966e-11
+WAIGSD = -1.1447549e-10
+PAIGSD = 1.106978e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.16719143
+LKT1 = -9.8483841e-09
+WKT1 = -2.9771263e-08
+PKT1 = 4.6681341e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.408 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.34650766+dvth0p408_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-3.3770949e-10+dlvth0p408_hp'
+WVTH0 = '1.0711219e-08+dwvth0p408_hp'
+PVTH0 = '-1.0357749e-15+dpvth0p408_hp'
+K1 = '0.68554981*dk1factorp_hp'
+LK1 = '-3.2777685e-09*dk1factorp_hp'
+WK1 = '-2.6330608e-08*dk1factorp_hp'
+PK1 = '1.5536623e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.12037461
+LVOFF = -2.5228885e-09
+WVOFF = -4.1055118e-10
+NFACTOR = 0.6446555
+ETA0 = 0.66179053
+LETA0 = -3.2956473e-08
+WETA0 = -7.9084044e-08
+PETA0 = 7.250424e-15
+ETAB = -0.15
+U0 = '(0.006325734*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.883227e-10*du0factorp_hp'
+WU0 = '3.4633852e-10*du0factorp_hp'
+PU0 = '-4.1430994e-17*du0factorp_hp'
+UA = 4.6674571e-19
+LUA = -7.2309561e-27
+WUA = -3.534429e-26
+PUA = 1.0357749e-33
+UB = 1e-19
+UC = -1.3204816e-19
+LUC = -2.185179e-27
+WUC = 5.7108284e-27
+PUC = 1.0357749e-33
+EU = 2
+VSAT = '213505.31*dvsatfactorp_hp'
+LVSAT = '-0.0026917433*dvsatfactorp_hp'
+WVSAT = '0.0074083653*dvsatfactorp_hp'
+PVSAT = '-5.1788743e-10*dvsatfactorp_hp'
+A0 = 0.48212166
+LA0 = 1.2614443e-07
+WA0 = -4.1055118e-08
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.16341085
+LKETA = 1.883227e-08
+WKETA = 4.6950387e-08
+PKETA = -4.1430994e-15
+DWG = 0
+DWB = 0
+PCLM = 3.4081334
+LPCLM = -1.6647091e-07
+WPCLM = -3.6239168e-07
+PPCLM = 3.1073246e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.005687904
+LAIGSD = 2.2786173e-11
+WAIGSD = 1.6811312e-10
+PAIGSD = -1.0800646e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.29779252
+LKT1 = 6.5555371e-09
+WKT1 = 3.2133657e-08
+PKT1 = -3.1073246e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.508 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.28776838+dvth0p508_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-9.2100629e-09+dlvth0p508_hp'
+WVTH0 = '-2.2114227e-09+dwvth0p508_hp'
+PVTH0 = '9.1614289e-16+dpvth0p508_hp'
+K1 = '0.60210432*dk1factorp_hp'
+LK1 = '5.8664757e-09*dk1factorp_hp'
+WK1 = '-7.9726019e-09*dk1factorp_hp'
+PK1 = '-4.5807145e-16*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1221666
+LVOFF = -4.6050315e-09
+WVOFF = -1.6313774e-11
+PVOFF = 4.5807145e-16
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0077349398*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.6313253e-11*du0factorp_hp'
+UA = 4.3168394e-19
+LUA = -6.6871744e-27
+WUA = -2.76307e-26
+PUA = 9.1614289e-34
+UB = 1e-19
+UC = -1.4915382e-19
+LUC = 6.6871744e-27
+WUC = 9.4740733e-27
+PUC = -9.1614289e-34
+EU = 2
+VSAT = '288444.76*dvsatfactorp_hp'
+LVSAT = '-0.005045777*dvsatfactorp_hp'
+WVSAT = '-0.0090783133*dvsatfactorp_hp'
+A0 = 0.23096646
+LA0 = 8.4501567e-08
+WA0 = 1.4199026e-08
+PA0 = 9.1614289e-15
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.29187779
+LKETA = -2.4985715e-08
+WKETA = -5.3213115e-08
+PKETA = 5.4968573e-15
+DWG = 0
+DWB = 0
+PCLM = 1.495319
+LPCLM = 1.6413973e-08
+WPCLM = 5.842748e-08
+PPCLM = -9.1614289e-15
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0078181388
+LAIGC = 3.3314287e-11
+WAIGC = -1.4990546e-11
+PAIGC = -7.3291431e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0075123204
+LAIGSD = -1.7074551e-10
+WAIGSD = -2.3325849e-10
+PAIGSD = 3.1776325e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.072056612
+LKT1 = -2.0061523e-08
+WKT1 = -1.7528244e-08
+PKT1 = 2.7484287e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.82080809
+LUTE = -1.2492858e-08
+WUTE = -2.842222e-08
+PUTE = 2.7484287e-15
+UA1 = 0
+UB1 = -1e-18
+UC1 = 4e-28
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.608 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.35359268+dvth0p608_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '8.779652e-09+dlvth0p608_hp'
+WVTH0 = '6.8065065e-09+dwvth0p608_hp'
+PVTH0 = '-1.5484481e-15+dpvth0p608_hp'
+K1 = '0.77767521*dk1factorp_hp'
+LK1 = '-2.0082193e-08*dk1factorp_hp'
+WK1 = '-3.2025813e-08*dk1factorp_hp'
+PK1 = '3.0968961e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.19220573
+LVOFF = 9.7020201e-09
+WVOFF = 9.5790473e-09
+PVOFF = -1.5019946e-15
+NFACTOR = 0.6446555
+ETA0 = 0.15815254
+LETA0 = 2.2605081e-08
+WETA0 = 1.9750613e-08
+PETA0 = -3.0968961e-15
+ETAB = -0.15
+U0 = '(0.017370729*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.4693303e-09*du0factorp_hp'
+WU0 = '-1.2837898e-09*du0factorp_hp'
+PU0 = '2.0129825e-16*du0factorp_hp'
+UA = -2.3356759e-18
+LUA = 3.3907622e-25
+WUA = 3.5149759e-25
+PUA = -4.6453442e-32
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '294262.23*dvsatfactorp_hp'
+LVSAT = '-0.016348318*dvsatfactorp_hp'
+WVSAT = '-0.0098753065*dvsatfactorp_hp'
+PVSAT = '1.5484481e-09*dvsatfactorp_hp'
+A0 = -1.1070416
+LA0 = 3.7742412e-07
+WA0 = 1.9750613e-07
+PA0 = -3.0968961e-14
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.28139101
+LKETA = -3.0072831e-08
+WKETA = -5.1776426e-08
+PKETA = 6.1937922e-15
+DWG = 0
+DWB = 0
+PCLM = 3.3634476
+LPCLM = -2.7650858e-07
+WPCLM = -1.9750613e-07
+PPCLM = 3.0968961e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0069878935
+LAIGC = 9.2842298e-11
+WAIGC = 9.8753065e-11
+PAIGC = -1.5484481e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0029744491
+LAIGSD = 3.3536758e-10
+WAIGSD = 3.8842988e-10
+PAIGSD = -3.7561169e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = 0.16041265
+LKT1 = -5.6512703e-08
+WKT1 = -4.9376532e-08
+PKT1 = 7.7422403e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.91138702
+LUTE = -3.733875e-09
+WUTE = -1.6012906e-08
+PUTE = 1.5484481e-15
+UA1 = 0
+UB1 = -1e-18
+UC1 = 7.2082529e-19
+LUC1 = -1.1302541e-25
+WUC1 = -9.8753064e-26
+PUC1 = 1.5484481e-32
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.708 PMOS
+LMIN = '1.38700000e-07+dlminp_hp'
+LMAX = '1.98800000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.2928203+dvth0p708_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.045777e-09+dlvth0p708_hp'
+K1 = '0.49173045*dk1factorp_hp'
+LK1 = '7.5686656e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.10667852
+LVOFF = -3.7086461e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3344973
+LETA0 = -5.045777e-09
+ETAB = -0.15
+U0 = '(0.0059083195*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.2797551e-10*du0factorp_hp'
+UA = 8.0269551e-19
+LUA = -7.5686656e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '206089.85*dvsatfactorp_hp'
+LVSAT = '-0.0025228885*dvsatfactorp_hp'
+A0 = 0.65640599
+LA0 = 1.0091554e-07
+AGS = -0.14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.1808985
+LKETA = 2.5228885e-08
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0078696173
+LAIGC = -4.5411993e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006442573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.28044925
+LKT1 = 1.2614443e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -1.0543594
+LUTE = 1.0091554e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = -1.608985e-19
+LUC1 = 2.5228885e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p708_hp'
+PVTH0 = '0.0+dpvth0p708_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.009 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32697544+dvth0p009_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.0422518e-09+dlvth0p009_hp'
+K1 = '0.63395087*dk1factorp_hp'
+LK1 = '4.0845036e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1273306
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0088722108*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.8380266e-10*du0factorp_hp'
+UA = 3.4e-19
+UB = 1e-19
+UC = -1.4604913e-19
+LUC = 4.0845036e-27
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.8395087
+LA0 = 4.0845036e-08
+AGS = -0.05185261
+LAGS = -1.2253511e-08
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.01604913
+LKETA = 4.0845036e-09
+DWG = 0
+DWB = 0
+PCLM = 2.5209826
+LPCLM = -8.1690072e-08
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.20395087
+LKT1 = -4.0845036e-09
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p009_hp'
+PVTH0 = '0.0+dpvth0p009_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.109 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.33250422+dvth0p109_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.1753379e-09+dlvth0p109_hp'
+WVTH0 = '5.512201e-08+dwvth0p109_hp'
+PVTH0 = '-8.6431311e-15+dpvth0p109_hp'
+K1 = '0.63395087*dk1factorp_hp'
+LK1 = '4.0845036e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1350709
+LVOFF = 1.2136794e-09
+WVOFF = 7.7170814e-08
+PVOFF = -1.2100384e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0090380745*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.0981008e-10*du0factorp_hp'
+WU0 = '-1.6536603e-09*du0factorp_hp'
+PU0 = '2.5929393e-16*du0factorp_hp'
+UA = 3.4e-19
+UB = 1e-19
+UC = -1.4604913e-19
+LUC = 4.0845036e-27
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.8395087
+LA0 = 4.0845036e-08
+AGS = -0.045039927
+LAGS = -1.3987338e-08
+WAGS = -6.7922445e-08
+PAGS = 1.7286262e-14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.01604913
+LKETA = 4.0845036e-09
+DWG = 0
+DWB = 0
+PCLM = 2.4528558
+LPCLM = -6.4351795e-08
+WPCLM = 6.7922445e-07
+PPCLM = -1.7286262e-13
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0061219589
+LAIGSD = -1.5604449e-11
+WAIGSD = -7.9147764e-10
+PAIGSD = 1.5557636e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.1928933
+LKT1 = -5.8183313e-09
+WKT1 = -1.1024402e-07
+PKT1 = 1.7286262e-14
+KT1L = 0
+KT2 = -0.04
+UTE = -0.92956195
+LUTE = -5.2014831e-09
+WUTE = -2.0376734e-07
+PUTE = 5.1858787e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.209 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31395087+dvth0p209_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-4.0845036e-09+dlvth0p209_hp'
+K1 = '0.62614709*dk1factorp_hp'
+LK1 = '6.0705654e-09*dk1factorp_hp'
+WK1 = '2.3185028e-08*dk1factorp_hp'
+PK1 = '-5.9005895e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.097312403
+LVOFF = -4.2493957e-09
+WVOFF = -3.5009687e-08
+PVOFF = 4.1304127e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0088614602*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.8211696e-10*du0factorp_hp'
+WU0 = '-1.1289393e-09*du0factorp_hp'
+PU0 = '1.7701769e-16*du0factorp_hp'
+UA = 3.4e-19
+UB = 1e-19
+UC = -1.5871534e-19
+LUC = 6.0705654e-27
+WUC = 3.7631311e-26
+PUC = -5.9005895e-33
+EU = 2
+VSAT = '207196.22*dvsatfactorp_hp'
+LVSAT = '0.0019860618*dvsatfactorp_hp'
+WVSAT = '0.023185028*dvsatfactorp_hp'
+PVSAT = '-5.9005895e-09*dvsatfactorp_hp'
+A0 = 0.99558428
+LA0 = 1.1238004e-09
+WA0 = -4.6370055e-07
+PA0 = 1.1801179e-13
+AGS = -0.083509298
+LAGS = -4.1968836e-09
+WAGS = 4.6370055e-08
+PAGS = -1.1801179e-14
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.01604913
+LKETA = 4.0845036e-09
+DWG = 0
+DWB = 0
+PCLM = 2.6814739
+LPCLM = -1.2253511e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0059282961
+LAIGSD = 2.5355175e-11
+WAIGSD = -2.1610533e-10
+PAIGSD = 3.3885315e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23
+KT1L = 0
+KT2 = -0.04
+UTE = -1.0215587
+LUTE = 1.8211696e-08
+WUTE = 6.9555083e-08
+PUTE = -1.7701769e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p209_hp'
+PVTH0 = '0.0+dpvth0p209_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.309 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32634775+dvth0p309_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.1406736e-09+dlvth0p309_hp'
+WVTH0 = '1.2049763e-08+dwvth0p309_hp'
+PVTH0 = '-1.8894028e-15+dpvth0p309_hp'
+K1 = '0.66903614*dk1factorp_hp'
+WK1 = '-1.8503133e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.13448212
+LVOFF = 7.7753201e-10
+WVOFF = 1.1192785e-09
+PVOFF = -7.5576111e-16
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0077*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 3.4575761e-19
+LUA = -3.88766e-27
+WUA = -5.5963927e-27
+PUA = 3.7788056e-33
+UB = 1e-19
+UC = -1.2e-19
+EU = 2
+VSAT = '231049.13*dvsatfactorp_hp'
+LVSAT = '-0.0040845036*dvsatfactorp_hp'
+A0 = 0.36576932
+LA0 = 1.6141171e-07
+WA0 = 1.4847959e-07
+PA0 = -3.7788056e-14
+AGS = -0.03580348
+LAGS = -1.6338014e-08
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.031324808
+LKETA = 7.9721636e-09
+WKETA = 1.4847959e-08
+PKETA = -3.7788056e-15
+DWG = 0
+DWB = 0
+PCLM = 2.8342307
+LPCLM = -1.6141171e-07
+WPCLM = -1.4847959e-07
+PPCLM = 3.7788056e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.00538558
+LAIGSD = 1.1753122e-10
+WAIGSD = 3.1141467e-10
+PAIGSD = -5.5709797e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2795875
+LKT1 = 7.7753201e-09
+WKT1 = 4.819905e-08
+PKT1 = -7.5576111e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.409 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.28702548+dvth0p409_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-9.6645144e-09+dlvth0p409_hp'
+WVTH0 = '-6.5889893e-09+dwvth0p409_hp'
+PVTH0 = '1.6768978e-15+dpvth0p409_hp'
+K1 = '0.68720791*dk1factorp_hp'
+LK1 = '-3.537759e-09*dk1factorp_hp'
+WK1 = '-2.7116548e-08*dk1factorp_hp'
+PK1 = '1.6768978e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.14479198
+LVOFF = 1.3057547e-09
+WVOFF = 6.0061495e-09
+PVOFF = -1.0061387e-15
+NFACTOR = 0.6446555
+ETA0 = 0.45160894
+WETA0 = -3.2844094e-08
+ETAB = -0.15
+U0 = '(0.0073011493*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.537759e-11*du0factorp_hp'
+WU0 = '1.8905525e-10*du0factorp_hp'
+PU0 = '-1.6768978e-17*du0factorp_hp'
+UA = 3.4945631e-19
+LUA = 1.1160022e-26
+WUA = -7.3495805e-27
+PUA = -3.3537955e-33
+UB = 1e-19
+UC = -1.4598425e-19
+WUC = 1.2316535e-26
+EU = 2
+VSAT = '244949.95*dvsatfactorp_hp'
+LVSAT = '-0.0076222626*dvsatfactorp_hp'
+WVSAT = '-0.0065889893*dvsatfactorp_hp'
+PVSAT = '1.6768978e-09*dvsatfactorp_hp'
+A0 = 0.54000919
+LA0 = 1.1706766e-07
+WA0 = 6.5889893e-08
+PA0 = -1.6768978e-14
+AGS = -0.013241241
+LAGS = -1.9875773e-08
+WAGS = -1.0694501e-08
+PAGS = 1.6768978e-15
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.080785226
+LKETA = -1.9457675e-08
+WKETA = -3.8292197e-08
+PKETA = 9.2229377e-15
+DWG = 0
+DWB = 0
+PCLM = 3.3186841
+LPCLM = -1.5244525e-07
+WPCLM = -3.7811049e-07
+PPCLM = 3.3537955e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.00637856
+LAIGSD = -8.5508697e-11
+WAIGSD = -1.5925785e-10
+PAIGSD = 4.0531122e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.13619928
+LKT1 = -1.8782284e-08
+WKT1 = -1.9766968e-08
+PKT1 = 5.0306933e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.90487552
+LUTE = -7.075518e-09
+WUTE = -2.1389002e-08
+PUTE = 3.3537955e-15
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.509 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31198308+dvth0p509_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.4131975e-09+dlvth0p509_hp'
+WVTH0 = '-1.0983179e-09+dwvth0p509_hp'
+PVTH0 = '7.4160806e-16+dpvth0p509_hp'
+K1 = '0.57047219*dk1factorp_hp'
+LK1 = '1.0826395e-08*dk1factorp_hp'
+WK1 = '-1.4346894e-09*dk1factorp_hp'
+PK1 = '-1.4832161e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.09629871
+LVOFF = -8.661116e-09
+WVOFF = -4.6623689e-09
+PVOFF = 1.1865729e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0071354959*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '9.3992793e-11*du0factorp_hp'
+WU0 = '2.2549898e-10*du0factorp_hp'
+PU0 = '-2.9664322e-17*du0factorp_hp'
+UA = 4.5808203e-19
+LUA = -1.0826395e-26
+WUA = -3.1247238e-26
+PUA = 1.4832161e-33
+UB = 1e-19
+UC = -1.0650602e-19
+WUC = 3.6313253e-27
+EU = 2
+VSAT = '213268.3*dvsatfactorp_hp'
+LVSAT = '0.0067418915*dvsatfactorp_hp'
+WVSAT = '0.00038097323*dvsatfactorp_hp'
+PVSAT = '-1.4832161e-09*dvsatfactorp_hp'
+A0 = 1.3693234
+LA0 = -9.3992793e-08
+WA0 = -1.1655922e-07
+PA0 = 2.9664322e-14
+AGS = -0.018855853
+LAGS = -1.8995402e-08
+WAGS = -9.4592865e-09
+PAGS = 1.4832161e-15
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.21712453
+LKETA = 5.4825849e-08
+WKETA = 2.7247949e-08
+PKETA = -7.1194374e-15
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0079446089
+LAIGC = 1.3483783e-11
+WAIGC = -4.2813957e-11
+PAIGC = -2.9664322e-18
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0050014398
+LAIGSD = 2.2296056e-10
+WAIGSD = 1.4370859e-10
+PAIGSD = -2.7332113e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.26904589
+LKT1 = 1.0826395e-08
+WKT1 = 9.4592865e-09
+PKT1 = -1.4832161e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.95258019
+LUTE = 8.1690072e-09
+WUTE = -1.0893976e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.609 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.35595005+dvth0p609_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '9.149288e-09+dlvth0p609_hp'
+WVTH0 = '4.925157e-09+dwvth0p609_hp'
+PVTH0 = '-1.2534525e-15+dpvth0p609_hp'
+K1 = '0.6496*dk1factorp_hp'
+WK1 = '-1.22752e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1303306
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0087814739*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.2253511e-10*du0factorp_hp'
+UA = 8.7710092e-19
+LUA = -1.6468718e-25
+WUA = -8.8652826e-26
+PUA = 2.2562144e-32
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '216049.13*dvsatfactorp_hp'
+LVSAT = '-0.0040845036*dvsatfactorp_hp'
+A0 = 0.5185261
+LA0 = 1.2253511e-07
+AGS = -0.08790174
+LAGS = -8.1690072e-09
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.010324463
+LKETA = 1.5668156e-08
+WKETA = -1.0836602e-09
+PKETA = -1.7548334e-15
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0087990993
+LAIGC = -1.9115477e-10
+WAIGC = -1.5987914e-10
+PAIGC = 2.5069049e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0012893312
+LAIGSD = 5.9959407e-10
+WAIGSD = 6.5226747e-10
+PAIGSD = -7.8930904e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2
+KT1L = 0
+KT2 = -0.04
+UTE = 0.063002661
+LUTE = -1.5651818e-07
+WUTE = -1.5002883e-07
+PUTE = 2.2562144e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.709 PMOS
+LMIN = '1.98800000e-07+dlminp_hp'
+LMAX = '2.96500000e-07+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31197544+dvth0p709_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.0422518e-09+dlvth0p709_hp'
+K1 = '0.54*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1303306
+NFACTOR = 0.6446555
+ETA0 = 0.3023176
+ETAB = -0.15
+U0 = '(0.0087814739*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.2253511e-10*du0factorp_hp'
+UA = 8.555783e-20
+LUA = 3.6760532e-26
+UB = 1e-19
+UC = -8e-20
+EU = 2
+VSAT = '216049.13*dvsatfactorp_hp'
+LVSAT = '-0.0040845036*dvsatfactorp_hp'
+A0 = 0.5185261
+LA0 = 1.2253511e-07
+AGS = -0.08790174
+LAGS = -8.1690072e-09
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.02
+DWG = 0
+DWB = 0
+PCLM = 1.6
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.007371607
+LAIGC = 3.2676029e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0071131479
+LAIGSD = -1.0514615e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2
+KT1L = 0
+KT2 = -0.04
+UTE = -1.2765404
+LUTE = 4.4929539e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 2.6049129e-20
+LUC1 = -4.0845034e-27
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p709_hp'
+PVTH0 = '0.0+dpvth0p709_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.010 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31457356+dvth0p010_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.1985288e-09+dlvth0p010_hp'
+K1 = '0.63638237*dk1factorp_hp'
+LK1 = '3.4656859e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.097371822
+LVOFF = -7.6245089e-09
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0082180881*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.7328429e-11*du0factorp_hp'
+UA = 3.4e-19
+UB = 1e-19
+UC = -2.2532338e-19
+LUC = 2.4259801e-26
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.65955935
+LA0 = 8.6642146e-08
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.027235252
+LKETA = -6.9313717e-09
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0057122462
+LAIGSD = 8.4068182e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.22
+KT1L = 0
+KT2 = -0.04
+UTE = -1.0180881
+LUTE = 1.7328429e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p010_hp'
+PVTH0 = '0.0+dpvth0p010_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.110 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31380574+dvth0p110_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.9341019e-09+dlvth0p110_hp'
+WVTH0 = '-7.6551817e-09+dwvth0p110_hp'
+PVTH0 = '7.3336641e-15+dpvth0p110_hp'
+K1 = '0.63638237*dk1factorp_hp'
+LK1 = '3.4656859e-09*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.093406604
+LVOFF = -9.3898844e-09
+WVOFF = -3.9533223e-08
+PVOFF = 1.7600794e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0082817615*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.7328429e-11*du0factorp_hp'
+WU0 = '-6.3482362e-10*du0factorp_hp'
+PU0 = '2.5443759e-30*du0factorp_hp'
+UA = 3.4e-19
+UB = 1e-19
+UC = -2.7156767e-19
+LUC = 3.6028971e-26
+WUC = 4.610555e-25
+PUC = -1.1733863e-31
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.65955935
+LA0 = 8.6642146e-08
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.027235252
+LKETA = -6.9313717e-09
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0056768058
+LAIGSD = 9.7687024e-11
+WAIGSD = 3.533405e-10
+PAIGSD = -1.3577986e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.22731618
+LKT1 = 2.9422925e-09
+WKT1 = 7.2942301e-08
+PKT1 = -2.9334656e-14
+KT1L = 0
+KT2 = -0.042890268
+LKT2 = 7.3557313e-10
+WKT2 = 2.8815969e-08
+PKT2 = -7.3336641e-15
+UTE = -1.0180881
+LUTE = 1.7328429e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.210 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31969311+dvth0p210_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.6231029e-09+dlvth0p210_hp'
+WVTH0 = '9.8362042e-09+dwvth0p210_hp'
+PVTH0 = '-2.503314e-15+dpvth0p210_hp'
+K1 = '0.6297609*dk1factorp_hp'
+LK1 = '5.1508518e-09*dk1factorp_hp'
+WK1 = '1.9672408e-08*dk1factorp_hp'
+PK1 = '-5.0066279e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.10237826
+LVOFF = -2.9601361e-09
+WVOFF = -1.2878446e-08
+PVOFF = -1.5019884e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0082470685*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.5754259e-11*du0factorp_hp'
+WU0 = '-5.3175054e-10*du0factorp_hp'
+PU0 = '2.503314e-17*du0factorp_hp'
+UA = 3.4e-19
+UB = 1e-19
+UC = -1.1462333e-19
+LUC = -5.1508518e-27
+WUC = -5.2261252e-27
+PUC = 5.0066279e-33
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.65955935
+LA0 = 8.6642146e-08
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.040478206
+LKETA = -1.0301704e-08
+WKETA = -3.9344817e-08
+PKETA = 1.0013256e-14
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0057525265
+LAIGSD = 7.008852e-11
+WAIGSD = 1.2837411e-10
+PAIGSD = -5.3784702e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.20938622
+LKT1 = -5.2462058e-09
+WKT1 = 1.9672408e-08
+PKT1 = -5.0066279e-15
+KT1L = 0
+KT2 = -0.029880448
+LKT2 = -2.5754259e-09
+WKT2 = -9.8362042e-09
+PKT2 = 2.503314e-15
+UTE = -1.0313311
+LUTE = 2.0698761e-08
+WUTE = 3.9344817e-08
+PUTE = -1.0013256e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.310 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.3143326+dvth0p310_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-5.1985288e-09+dlvth0p310_hp'
+WVTH0 = '4.6257831e-09+dwvth0p310_hp'
+K1 = '0.66255547*dk1factorp_hp'
+LK1 = '1.6493324e-09*dk1factorp_hp'
+WK1 = '-1.2203914e-08*dk1factorp_hp'
+PK1 = '-1.6031511e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1292777
+LVOFF = -5.4699379e-10
+WVOFF = 1.3267811e-08
+PVOFF = -3.8475627e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0075703864*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '3.2986649e-11*du0factorp_hp'
+WU0 = '1.2598437e-10*du0factorp_hp'
+PU0 = '-3.2063022e-17*du0factorp_hp'
+UA = 3.3696261e-19
+LUA = -1.6493324e-27
+WUA = 2.9523477e-27
+PUA = 1.6031511e-33
+UB = 1e-19
+UC = -1.2e-19
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.65955935
+LA0 = 8.6642146e-08
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0057342376
+LAIGSD = 2.879787e-11
+WAIGSD = 1.4615099e-10
+PAIGSD = -1.3650191e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.1692992
+LKT1 = -2.0293052e-08
+WKT1 = -1.9292179e-08
+PKT1 = 9.6189067e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.90012339
+LUTE = -1.2693596e-08
+WUTE = -8.818906e-08
+PUTE = 2.2444116e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+PVTH0 = '0.0+dpvth0p310_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.410 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31636836+dvth0p410_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-2.1967536e-09+dlvth0p410_hp'
+WVTH0 = '5.5907325e-09+dwvth0p410_hp'
+PVTH0 = '-1.4228414e-15+dpvth0p410_hp'
+K1 = '0.6742185*dk1factorp_hp'
+LK1 = '-2.3195535e-10*dk1factorp_hp'
+WK1 = '-1.7732193e-08*dk1factorp_hp'
+PK1 = '-7.1142071e-16*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.10561724
+LVOFF = -8.6642146e-09
+WVOFF = 2.0527559e-09
+NFACTOR = 0.6446555
+ETA0 = 0.35725058
+LETA0 = 2.4014201e-08
+WETA0 = 1.1881766e-08
+PETA0 = -1.1382731e-14
+ETAB = -0.15
+U0 = '(0.006986594*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.154319e-10*du0factorp_hp'
+WU0 = '4.0270198e-10*du0factorp_hp'
+PU0 = '-7.1142071e-17*du0factorp_hp'
+UA = 3.275243e-19
+LUA = 1.6741719e-26
+WUA = 7.4261035e-27
+PUA = -7.1142071e-33
+UB = 1e-19
+UC = -1.1059987e-19
+LUC = -9.0053255e-27
+WUC = -4.4556621e-27
+PUC = 4.2685243e-33
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.65955935
+LA0 = 8.6642146e-08
+AGS = -0.10313338
+LAGS = 3.0017752e-09
+WAGS = 1.4852207e-09
+PAGS = -1.4228414e-15
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.0015666885
+LKETA = 1.5008876e-09
+WKETA = 7.4261035e-10
+PKETA = -7.1142071e-16
+DWG = 0
+DWB = 0
+PCLM = 2.0119974
+LPCLM = 1.8010651e-07
+WPCLM = 8.9113241e-08
+PPCLM = -8.5370485e-14
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006042573
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.22179479
+LKT1 = 3.0017752e-09
+WKT1 = 5.5907325e-09
+PKT1 = -1.4228414e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -1.033469
+LUTE = 2.5651533e-08
+WUTE = -2.4983221e-08
+PUTE = 4.2685243e-15
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.510 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.2879703+dvth0p510_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.1524449e-08+dlvth0p510_hp'
+WVTH0 = '-6.5683887e-10+dwvth0p510_hp'
+PVTH0 = '6.2925164e-16+dpvth0p510_hp'
+K1 = '0.71653882*dk1factorp_hp'
+LK1 = '-2.6347564e-08*dk1factorp_hp'
+WK1 = '-2.7042663e-08*dk1factorp_hp'
+PK1 = '5.0340131e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.096286535
+LVOFF = -8.6642146e-09
+NFACTOR = 0.6446555
+ETA0 = 0.41125861
+LETA0 = -2.7725487e-08
+ETAB = -0.15
+U0 = '(0.008097104*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.5073646e-10*du0factorp_hp'
+WU0 = '1.5838979e-10*du0factorp_hp'
+PU0 = '-1.2585033e-17*du0factorp_hp'
+UA = 3.5319641e-19
+LUA = 1.5866995e-26
+WUA = 1.7782396e-27
+PUA = -6.921768e-33
+UB = 1e-19
+UC = -1.2488162e-19
+LUC = 4.6765881e-27
+WUC = -1.3136777e-27
+PUC = 1.2585033e-33
+EU = 2
+VSAT = '206043.11*dvsatfactorp_hp'
+LVSAT = '0.0085807041*dvsatfactorp_hp'
+WVSAT = '0.0019705166*dvsatfactorp_hp'
+PVSAT = '-1.8877549e-09*dvsatfactorp_hp'
+A0 = 0.70451392
+LA0 = 7.5201208e-08
+WA0 = -9.8900061e-09
+PA0 = 2.5170065e-15
+AGS = -0.10235364
+LAGS = 2.2547836e-09
+WAGS = 1.3136777e-09
+PAGS = -1.2585033e-15
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.00061456059
+LKETA = -5.8874904e-10
+WKETA = 2.6273555e-10
+PKETA = -2.5170065e-16
+DWG = 0
+DWB = 0
+PCLM = 2.4170576
+LPCLM = -2.0794115e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076604311
+LAIGC = 8.5807041e-11
+WAIGC = 1.9705166e-11
+PAIGC = -1.8877549e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0061022856
+LAIGSD = -5.7204694e-11
+WAIGSD = -1.3136777e-11
+PAIGSD = 1.2585033e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.19041111
+LKT1 = -9.1861553e-09
+WKT1 = -1.3136777e-09
+PKT1 = 1.2585033e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -1.0525565
+LUTE = 3.3612977e-08
+WUTE = -2.0783982e-08
+PUTE = 2.5170065e-15
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.610 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.29276475+dvth0p610_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-6.9313717e-09+dlvth0p610_hp'
+K1 = '0.60874712*dk1factorp_hp'
+LK1 = '1.0397058e-08*dk1factorp_hp'
+WK1 = '-1.22752e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = 0.013526003
+LVOFF = -3.6611505e-08
+WVOFF = -1.5044318e-08
+PVOFF = 3.8287788e-15
+NFACTOR = 1.498753
+LNFACTOR = -2.1736782e-07
+WNFACTOR = -1.1701136e-07
+PNFACTOR = 2.9779391e-14
+ETA0 = 0.41125861
+LETA0 = -2.7725487e-08
+ETAB = -0.15
+U0 = '(0.0086431642*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-8.7335284e-11*du0factorp_hp'
+WU0 = '8.3579542e-11*du0factorp_hp'
+PU0 = '-2.1270994e-17*du0factorp_hp'
+UA = 5.4919716e-19
+LUA = -8.1235676e-26
+WUA = -2.5073863e-26
+PUA = 6.3812981e-33
+UB = 1e-19
+UC = -1.344705e-19
+LUC = 1.3862743e-26
+EU = 2
+VSAT = '220426.44*dvsatfactorp_hp'
+LVSAT = '-0.0051985288*dvsatfactorp_hp'
+A0 = 0.63232409
+LA0 = 9.3573518e-08
+AGS = -0.092764748
+LAGS = -6.9313717e-09
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = -0.018536716
+LKETA = 1.7758174e-08
+WKETA = 2.8864605e-09
+PKETA = -2.7652292e-15
+DWG = 0
+DWB = 0
+PCLM = 2.4170576
+LPCLM = -2.0794115e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0076421947
+LAIGC = 1.0327744e-10
+WAIGC = 2.2203542e-11
+PAIGC = -2.1270994e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0077796113
+LAIGSD = -1.0521822e-09
+WAIGSD = -2.429304e-10
+PAIGSD = 1.4889695e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.26100697
+LKT1 = 1.5526273e-08
+WKT1 = 8.3579542e-09
+PKT1 = -2.1270994e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -1.0612992
+LUTE = 1.2961665e-07
+WUTE = -1.9586229e-08
+PUTE = -1.0635497e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p610_hp'
+PVTH0 = '0.0+dpvth0p610_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.710 PMOS
+LMIN = '2.96500000e-07+dlminp_hp'
+LMAX = '1.00000000e-06+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.29276475+dvth0p710_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-6.9313717e-09+dlvth0p710_hp'
+K1 = '0.49914712*dk1factorp_hp'
+LK1 = '1.0397058e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.12079826
+LVOFF = -2.4259801e-09
+NFACTOR = 0.45400873
+LNFACTOR = 4.8519602e-08
+ETA0 = 0.41125861
+LETA0 = -2.7725487e-08
+ETAB = -0.15
+U0 = '(0.0093894101*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-2.7725487e-10*du0factorp_hp'
+UA = 3.2532338e-19
+LUA = -2.4259801e-26
+UB = 1e-19
+UC = -1.344705e-19
+LUC = 1.3862743e-26
+EU = 2
+VSAT = '220426.44*dvsatfactorp_hp'
+LVSAT = '-0.0051985288*dvsatfactorp_hp'
+A0 = 0.63232409
+LA0 = 9.3573518e-08
+AGS = -0.092764748
+LAGS = -6.9313717e-09
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.0072352523
+LKETA = -6.9313717e-09
+DWG = 0
+DWB = 0
+PCLM = 2.4170576
+LPCLM = -2.0794115e-07
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0078404407
+LAIGC = -8.6642146e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0056105899
+LAIGSD = 2.7725487e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.18638237
+LKT1 = -3.4656859e-09
+KT1L = 0
+KT2 = -0.04
+UTE = -1.2361763
+LUTE = 3.4656859e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1e-20
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p710_hp'
+PVTH0 = '0.0+dpvth0p710_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.011 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32+dvth0p011_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.62521*dk1factorp_hp'
+LK1 = '1.416882e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1201206
+LVOFF = 1.416882e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0083479*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.416882e-10*du0factorp_hp'
+UA = 4.2874e-19
+LUA = -8.501292e-26
+UB = 1e-19
+UC = -2e-19
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.03479
+LKETA = -1.416882e-08
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0058
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.20521
+LKT1 = -1.416882e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.94084
+LUTE = -5.667528e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.1353e-19
+LUC1 = -9.918174e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p011_hp'
+WVTH0 = '0.0+dwvth0p011_hp'
+PVTH0 = '0.0+dpvth0p011_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.111 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32+dvth0p111_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.62521*dk1factorp_hp'
+LK1 = '1.416882e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.12113725
+LVOFF = 1.7176076e-08
+WVOFF = 1.0136017e-08
+PVOFF = -2.9982339e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0084429644*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.7176076e-10*du0factorp_hp'
+WU0 = '-9.4779166e-10*du0factorp_hp'
+PU0 = '2.9982339e-16*du0factorp_hp'
+UA = 4.2874e-19
+LUA = -8.501292e-26
+UB = 1e-19
+UC = -1.8373357e-19
+LUC = -4.811609e-26
+WUC = -1.6217627e-25
+PUC = 4.7971742e-31
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.041068195
+LKETA = -2.0183331e-08
+WKETA = -6.2593609e-08
+PKETA = 5.9964677e-14
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0057473846
+LAIGSD = 3.0072556e-11
+WAIGSD = 5.2457592e-10
+PAIGSD = -2.9982339e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2031767
+LKT1 = -2.0183331e-08
+WKT1 = -2.0272034e-08
+PKT1 = 5.9964677e-14
+KT1L = 0
+KT2 = -0.045261544
+LKT2 = 3.0072556e-09
+WKT2 = 5.2457592e-08
+PKT2 = -2.9982339e-14
+UTE = -0.92828361
+LUTE = -6.8704302e-08
+WUTE = -1.2518722e-07
+PUTE = 1.1992935e-13
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.6375556e-19
+LUC1 = -1.4729783e-25
+WUC1 = -5.0074887e-25
+PUC1 = 4.7971741e-31
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p111_hp'
+WVTH0 = '0.0+dwvth0p111_hp'
+PVTH0 = '0.0+dpvth0p111_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.211 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32243122+dvth0p211_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '7.2231416e-09+dwvth0p211_hp'
+K1 = '0.6275391*dk1factorp_hp'
+LK1 = '7.2793287e-09*dk1factorp_hp'
+WK1 = '-6.9197696e-09*dk1factorp_hp'
+PK1 = '2.0468679e-14*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1200547
+LVOFF = 1.3973901e-08
+WVOFF = 6.9197696e-09
+PVOFF = -2.0468679e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0080424313*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.7028809e-10*du0factorp_hp'
+WU0 = '2.4219194e-10*du0factorp_hp'
+PU0 = '-7.1640375e-16*du0factorp_hp'
+UA = 4.2874e-19
+LUA = -8.501292e-26
+UB = 1e-19
+UC = -2.3832e-19
+LUC = 1.1335056e-25
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.73561693
+LA0 = 1.3778983e-08
+WA0 = 4.2732106e-08
+PA0 = -4.0937357e-14
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.015341791
+LKETA = 1.3778983e-08
+WKETA = 1.3839539e-08
+PKETA = -4.0937357e-14
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0058636802
+LAIGSD = -3.6396644e-11
+WAIGSD = 1.7906168e-10
+PAIGSD = -1.0234339e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2076709
+LKT1 = -6.8894913e-09
+WKT1 = -6.9197696e-09
+PKT1 = 2.0468679e-14
+KT1L = 0
+KT2 = -0.021578017
+LKT2 = -1.0529156e-08
+WKT2 = -1.7906168e-08
+PKT2 = 1.0234339e-14
+UTE = -0.96576179
+LUTE = -4.2116623e-08
+WUTE = -1.3839539e-08
+PUTE = 4.0937357e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = -4.7899994e-21
+LUC1 = 1.4168819e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p211_hp'
+PVTH0 = '0.0+dpvth0p211_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.311 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31975904+dvth0p311_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '4.6257831e-09+dwvth0p311_hp'
+K1 = '0.64103186*dk1factorp_hp'
+LK1 = '2.2268947e-08*dk1factorp_hp'
+WK1 = '-2.0034729e-08*dk1factorp_hp'
+PK1 = '5.89877e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.10837644
+LVOFF = -2.0570395e-08
+WVOFF = -4.4315002e-09
+PVOFF = 1.3108378e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0083371916*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-7.0161265e-10*du0factorp_hp'
+WU0 = '-4.4315002e-11*du0factorp_hp'
+PU0 = '1.3108378e-16*du0factorp_hp'
+UA = 4.3101958e-19
+LUA = -9.1755913e-26
+WUA = -2.2157501e-27
+PUA = 6.5541889e-33
+UB = 1e-19
+UC = -2.6647446e-19
+LUC = 1.4032253e-25
+WUC = 2.7366133e-26
+PUC = -2.6216755e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.80773446
+LA0 = -5.5309611e-08
+WA0 = -2.7366133e-08
+PA0 = 2.6216755e-14
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.02958
+LKETA = -2.833764e-08
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0061129013
+LAIGSD = -3.3396194e-10
+WAIGSD = -6.3181228e-11
+PAIGSD = 1.8689007e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.23342639
+LKT1 = 4.1140791e-08
+WKT1 = 1.8114567e-08
+PKT1 = -2.6216755e-14
+KT1L = 0
+KT2 = -0.04
+UTE = -0.98375964
+LUTE = 6.7429927e-08
+WUTE = 3.6543687e-09
+PUTE = -6.5541889e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = -6.1098915e-20
+LUC1 = 6.811276e-26
+WUC1 = 5.4732265e-26
+PUC1 = -5.243351e-32
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p311_hp'
+PVTH0 = '0.0+dpvth0p311_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.411 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31866142+dvth0p411_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '4.1055118e-09+dwvth0p411_hp'
+K1 = '0.61916604*dk1factorp_hp'
+LK1 = '5.2508308e-08*dk1factorp_hp'
+WK1 = '-9.6703278e-09*dk1factorp_hp'
+PK1 = '-8.4346874e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.11565119
+LVOFF = 9.4830685e-10
+WVOFF = -9.8327008e-10
+PVOFF = 2.9085129e-15
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.007678889*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-5.4778666e-10*du0factorp_hp'
+WU0 = '2.6772043e-10*du0factorp_hp'
+PU0 = '5.8170258e-17*du0factorp_hp'
+UA = 4.3915524e-19
+LUA = -9.0200716e-26
+WUA = -6.072052e-27
+PUA = 5.8170258e-33
+UB = 1e-19
+UC = -2.4717071e-19
+LUC = 1.2182954e-25
+WUC = 1.8216156e-26
+PUC = -1.7451077e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.02958
+LKETA = -2.833764e-08
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0059796075
+LAIGSD = 6.0320917e-11
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.20387142
+LKT1 = -1.416882e-08
+WKT1 = 4.1055118e-09
+PKT1 = -1.614549e-29
+KT1L = 0
+KT2 = -0.04
+UTE = -0.97117362
+LUTE = -3.4027481e-08
+WUTE = -2.3114031e-09
+PUTE = -1.7451077e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 5.437e-20
+LUC1 = -4.250646e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p411_hp'
+PVTH0 = '0.0+dpvth0p411_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.511 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.3+dvth0p511_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.62542133*dk1factorp_hp'
+LK1 = '6.0942997e-08*dk1factorp_hp'
+WK1 = '-1.1046492e-08*dk1factorp_hp'
+PK1 = '-1.0290319e-14*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1201206
+LVOFF = 1.416882e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0070149386*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.8597802e-10*du0factorp_hp'
+WU0 = '4.1378952e-10*du0factorp_hp'
+PU0 = '-2.5725797e-16*du0factorp_hp'
+UA = 5.2175747e-19
+LUA = -1.456145e-25
+WUA = -2.4244543e-26
+PUA = 1.8008058e-32
+UB = 1e-19
+UC = -2.1319482e-19
+LUC = 8.9280637e-26
+WUC = 1.074146e-26
+PUC = -1.0290319e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.73418723
+LA0 = 4.6774177e-08
+WA0 = 3.4788096e-09
+PA0 = -1.0290319e-14
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.02958
+LKETA = -2.833764e-08
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0062237316
+LAIGSD = -1.7354997e-10
+WAIGSD = -5.3707301e-11
+PAIGSD = 5.1451595e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.18521
+LKT1 = -1.416882e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -0.58178855
+LUTE = -4.1738271e-07
+WUTE = -8.7976118e-08
+PUTE = 6.6887073e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 5.437e-20
+LUC1 = -4.250646e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p511_hp'
+WVTH0 = '0.0+dwvth0p511_hp'
+PVTH0 = '0.0+dpvth0p511_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.611 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.2668704+dvth0p611_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-3.1738157e-08+dlvth0p611_hp'
+WVTH0 = '-4.5387552e-09+dwvth0p611_hp'
+PVTH0 = '4.3481275e-15+dpvth0p611_hp'
+K1 = '0.7006492*dk1factorp_hp'
+LK1 = '-7.7645134e-08*dk1factorp_hp'
+WK1 = '-2.135271e-08*dk1factorp_hp'
+PK1 = '8.696255e-15*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.05935836
+LVOFF = 3.3211714e-08
+WVOFF = -8.3244269e-09
+PVOFF = -2.6088765e-15
+NFACTOR = 1.2718555
+WNFACTOR = -8.59264e-08
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.010249892*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-1.6265805e-09*du0factorp_hp'
+WU0 = '-2.9399104e-11*du0factorp_hp'
+PU0 = '8.696255e-17*du0factorp_hp'
+UA = 2.804124e-19
+LUA = 1.7626012e-25
+WUA = 8.8197312e-27
+PUA = -2.6088765e-32
+UB = 1e-19
+UC = -3.335676e-19
+LUC = 2.0459776e-25
+WUC = 2.7232531e-26
+PUC = -2.6088765e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75958
+LA0 = -2.833764e-08
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.1620984
+LKETA = -1.5529027e-07
+WKETA = -1.8155021e-08
+PKETA = 1.739251e-14
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0042005733
+LAIGSD = 2.3765362e-09
+WAIGSD = 2.2346539e-10
+PAIGSD = -2.9791022e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.2962692
+LKT1 = 4.9307494e-08
+WKT1 = 1.521511e-08
+PKT1 = -8.696255e-15
+KT1L = 0
+KT2 = -0.04
+UTE = -0.99995
+LUTE = 7.08441e-08
+WUTE = -3.0688e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 5.437e-20
+LUC1 = -4.250646e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.711 PMOS
+LMIN = '1.00000000e-06+dlminp_hp'
+LMAX = '3.00000000e-06+dlmaxp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.307395+dvth0p711_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '7.08441e-09+dlvth0p711_hp'
+K1 = '0.51*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1336836
+LVOFF = 9.918174e-09
+NFACTOR = 0.5046555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0099874*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '-8.501292e-10*du0factorp_hp'
+UA = 3.5916e-19
+LUA = -5.667528e-26
+UB = 1e-19
+UC = -9.042e-20
+LUC = -2.833764e-26
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75958
+LA0 = -2.833764e-08
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0061958
+LAIGSD = -2.833764e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.16042
+LKT1 = -2.833764e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -1.27395
+LUTE = 7.08441e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 5.437e-20
+LUC1 = -4.250646e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+WVTH0 = '0.0+dwvth0p711_hp'
+PVTH0 = '0.0+dpvth0p711_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.012 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '1.00000000e-05+dwminp0_hp'
+WMAX = '1.01000000e-04+wmaxoffsetp_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32+dvth0p012_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.63*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1153306
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0080154857*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '8.4159326e-10*du0factorp_hp'
+UA = 4e-19
+UB = 1e-19
+UC = -1.0042e-19
+LUC = -2.9455764e-25
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.072677143
+LKETA = -1.2623899e-07
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077784514
+LAIGC = -8.4159326e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0058
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.21
+KT1L = 0
+KT2 = -0.04
+UTE = -0.98845143
+LUTE = 8.4159326e-08
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.0845143e-19
+LUC1 = -8.4159326e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p012_hp'
+WVTH0 = '0.0+dwvth0p012_hp'
+PVTH0 = '0.0+dpvth0p012_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.112 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '3.00000000e-06+dwminp1_hp'
+WMAX = '1.00000000e-05+dwmaxp1_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.32+dvth0p112_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.63*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.11231127
+LVOFF = -8.9311815e-09
+WVOFF = -3.0102731e-08
+PVOFF = 8.9043879e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0079796103*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+LU0 = '1.1988405e-09*du0factorp_hp'
+WU0 = '3.5767776e-10*du0factorp_hp'
+PU0 = '-3.5617552e-15*du0factorp_hp'
+UA = 3.8792268e-19
+LUA = 3.5724726e-26
+WUA = 1.2041093e-25
+PUA = -3.5617552e-31
+UB = 1e-19
+UC = -8.8342675e-20
+LUC = -3.3028237e-25
+WUC = -1.2041093e-25
+PUC = 3.5617552e-31
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.082960697
+LKETA = -1.4410135e-07
+WKETA = -1.0252704e-07
+PKETA = 1.7808776e-13
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077844901
+LAIGC = -1.0202169e-10
+WAIGC = -6.0205463e-11
+PAIGC = 1.7808776e-16
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0058179377
+LAIGSD = -1.7862363e-10
+WAIGSD = -1.7883888e-10
+PAIGSD = 1.7808776e-15
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.21
+KT1L = 0
+KT2 = -0.03820623
+LKT2 = -1.7862363e-08
+WKT2 = -1.7883888e-08
+PKT2 = 1.7808776e-13
+UTE = -1.010155
+LUTE = 1.7347114e-07
+WUTE = 2.1638416e-07
+PUTE = -8.9043879e-13
+UA1 = 0
+UB1 = -1e-18
+UC1 = 3.3714645e-20
+LUC1 = 2.3736321e-25
+WUC1 = 7.4512573e-25
+PUC1 = -3.2055796e-30
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p112_hp'
+WVTH0 = '0.0+dwvth0p112_hp'
+PVTH0 = '0.0+dpvth0p112_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.212 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '1.00000000e-06+dwminp2_hp'
+WMAX = '3.00000000e-06+dwmaxp2_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31897264+dvth0p212_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '-1.0230473e-08+dlvth0p212_hp'
+WVTH0 = '-3.0522933e-09+dwvth0p212_hp'
+PVTH0 = '3.0394736e-14+dpvth0p212_hp'
+K1 = '0.63*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.12244346
+LVOFF = 2.1039831e-08
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0081*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 4.2845143e-19
+LUA = -8.4159326e-26
+UB = 1e-19
+UC = -1.2195427e-19
+LUC = -2.3085926e-25
+WUC = -2.055087e-26
+PUC = 6.0789472e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75410945
+LA0 = -4.0921893e-08
+WA0 = -1.2209173e-08
+PA0 = 1.2157894e-13
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.06228574
+LKETA = -1.2508122e-07
+WKETA = -4.1101739e-08
+PKETA = 1.2157894e-13
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077573086
+LAIGC = -2.1618716e-11
+WAIGC = 2.055087e-11
+PAIGC = -6.0789472e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0057782901
+LAIGSD = 2.1618716e-10
+WAIGSD = -6.1045865e-11
+PAIGSD = 6.0789472e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.21
+KT1L = 0
+KT2 = -0.046280439
+LKT2 = 6.2540609e-08
+WKT2 = 6.1045865e-09
+PKT2 = -6.0789472e-14
+UTE = -0.90965423
+LUTE = -2.0808278e-07
+WUTE = -8.2203479e-08
+PUTE = 2.4315789e-13
+UA1 = 0
+UB1 = -1e-18
+UC1 = 3.6752015e-19
+LUC1 = -1.0871246e-24
+WUC1 = -2.4661044e-25
+PUC1 = 7.2947367e-31
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.312 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '5.00000000e-07+dwminp3_hp'
+WMAX = '1.00000000e-06+dwmaxp3_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.33364196+dvth0p312_hp+(mcm_PENHHP_vth0*mcmScale)'
+LVTH0 = '4.1065695e-08+dlvth0p312_hp'
+WVTH0 = '1.120629e-08+dwvth0p312_hp'
+PVTH0 = '-1.9465139e-14+dpvth0p312_hp'
+K1 = '0.64856024*dk1factorp_hp'
+WK1 = '-1.8040554e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.12921353
+LVOFF = 4.1065695e-08
+WVOFF = 6.5805069e-09
+PVOFF = -1.9465139e-14
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0081*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 4.4199157e-19
+LUA = -1.2421105e-25
+WUA = -1.3161014e-26
+PUA = 3.8930279e-32
+UB = 1e-19
+UC = -1.4859315e-19
+LUC = -2.0837038e-25
+WUC = 5.3421187e-27
+PUC = 3.8930279e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.66580375
+LA0 = 3.6452142e-07
+WA0 = 7.3623964e-08
+PA0 = -2.7251195e-13
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.0064598623
+LKETA = 4.0051727e-08
+WKETA = 1.3161014e-08
+PKETA = -3.8930279e-14
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0077784514
+LAIGC = -8.4159326e-11
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.005444683
+LAIGSD = 1.6426278e-09
+WAIGSD = 2.6322028e-10
+PAIGSD = -7.7860558e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.21951807
+WKT1 = 9.2515663e-09
+KT1L = 0
+KT2 = -0.04
+UTE = -0.98872971
+LUTE = 8.213139e-08
+WUTE = -5.3421187e-09
+PUTE = -3.8930279e-14
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.028137e-19
+LUC1 = -4.1674075e-25
+WUC1 = 1.0684238e-26
+PUC1 = 7.7860556e-32
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.412 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '2.40000000e-07+dwminp4_hp'
+WMAX = '5.00000000e-07+dwmaxp4_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.31866142+dvth0p412_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '4.1055118e-09+dwvth0p412_hp'
+K1 = '0.63691732*dk1factorp_hp'
+WK1 = '-1.2521811e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1153306
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0074937008*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '2.8738583e-10*du0factorp_hp'
+UA = 4.3520862e-19
+LUA = -7.8526615e-26
+WUA = -9.9458956e-27
+PUA = 1.7275855e-32
+UB = 1e-19
+UC = -1.5098562e-19
+LUC = -1.6268594e-25
+WUC = 6.4761516e-27
+PUC = 1.7275855e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.882736
+LA0 = -3.9263307e-07
+WA0 = -2.9201919e-08
+PA0 = 8.6379276e-14
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.046547199
+LKETA = -7.8526615e-08
+WKETA = -5.8403838e-09
+PKETA = 1.7275855e-14
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.0078030944
+LAIGC = -1.5705323e-10
+WAIGC = -1.1680768e-11
+PAIGC = 3.4551711e-17
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0059475437
+LAIGSD = 1.5516561e-10
+WAIGSD = 2.4864266e-11
+PAIGSD = -7.3548499e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.20866142
+WKT1 = 4.1055118e-09
+KT1L = 0
+KT2 = -0.04
+UTE = -0.88410529
+LUTE = -2.9157562e-07
+WUTE = -5.4934094e-08
+PUTE = 1.3820684e-13
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.2535429e-19
+LUC1 = -2.5247798e-25
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p412_hp'
+PVTH0 = '0.0+dpvth0p412_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.512 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '1.50000000e-07+dwminp5_hp'
+WMAX = '2.40000000e-07+dwmaxp5_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.3+dvth0p512_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.6460241*dk1factorp_hp'
+WK1 = '-1.4525301e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1153306
+NFACTOR = 0.6446555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0073144578*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+WU0 = '3.2681928e-10*du0factorp_hp'
+UA = 4.7253012e-19
+WUA = -1.8156627e-26
+UB = 1e-19
+UC = -1.3107962e-19
+LUC = -1.5361612e-25
+WUC = 2.096831e-27
+PUC = 1.5280494e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.02
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.006325589
+LAIGSD = -4.7484415e-10
+WAIGSD = -5.8305697e-11
+PAIGSD = 6.5053649e-17
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.213481
+LKT1 = 6.9456793e-08
+WKT1 = 5.1658196e-09
+PKT1 = -1.5280494e-14
+KT1L = 0
+KT2 = -0.04
+UTE = -1.2593552
+LUTE = 1.5868596e-06
+WUTE = 2.7620898e-08
+PUTE = -2.750489e-13
+UA1 = 0
+UB1 = -1e-18
+UC1 = 1.2535429e-19
+LUC1 = -2.5247798e-25
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p512_hp'
+WVTH0 = '0.0+dwvth0p512_hp'
+PVTH0 = '0.0+dpvth0p512_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.612 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '1.20000000e-07+dwminp6_hp'
+WMAX = '1.50000000e-07+dwmaxp6_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.2776+dvth0p612_hp+(mcm_PENHHP_vth0*mcmScale)'
+WVTH0 = '-3.0688e-09+dwvth0p612_hp'
+K1 = '0.6744*dk1factorp_hp'
+WK1 = '-1.84128e-08*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.0481306
+WVOFF = -9.2064e-09
+NFACTOR = 1.2718555
+WNFACTOR = -8.59264e-08
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0097*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 3.4e-19
+UB = 1e-19
+UC = -3.1390549e-19
+LUC = 1.4643723e-25
+WUC = 2.7143974e-26
+PUC = -2.5826814e-32
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0.1096
+WKETA = -1.22752e-08
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.004366688
+LAIGSD = 1.8851689e-09
+WAIGSD = 2.1006374e-10
+PAIGSD = -2.5826814e-16
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.13791189
+LKT1 = -4.1911344e-07
+WKT1 = -5.1871488e-09
+PKT1 = 5.1653628e-14
+KT1L = 0
+KT2 = -0.04
+UTE = -1.1523989
+LUTE = 5.2178782e-07
+WUTE = 1.2967872e-08
+PUTE = -1.2913407e-13
+UA1 = 0
+UB1 = -1e-18
+UC1 = 3.8027909e-19
+LUC1 = -1.0065455e-24
+WUC1 = -3.4924698e-26
+PUC1 = 1.0330726e-31
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p612_hp'
+PVTH0 = '0.0+dpvth0p612_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.MODEL PENHHP.712 PMOS
+LMIN = '3.00000000e-06+dlminp_hp'
+LMAX = '1.00000000e-05+lmaxoffsetp_hp'
+WMIN = '1.10000000e-07+wminoffsetp_hp'
+WMAX = '1.20000000e-07+dwmaxp7_hp'
+BINUNIT = 0
+LEVEL = 54
+VERSION = 4.5
+PARAMCHK = 0
+MOBMOD = 2
+CAPMOD = 2
+IGCMOD = 1
+IGBMOD = 1
+GEOMOD = 0
+DIOMOD = 1
+RDSMOD = 0
+RBODYMOD = 0
+RGATEMOD = 0
+PERMOD = 1
+ACNQSMOD = 0
+TRNQSMOD = 0
+TNOM = 23
+TOXE = '2.36e-09+dtoxp_hp'
+TOXP = '2.16e-09+dtoxp_hp'
+TOXM = 2.36e-09
+EPSROX = 3.9
+WINT = '1.49200000e-08+dwintp_hp'
+LINT = '2.10000000e-08+dlintp_hp'
+LL = 0
+WL = 0
+LLN = 1
+WLN = 1
+LW = 0
+WW = -9.454e-17
+LWN = 1
+WWN = 1.165
+LWL = 0
+WWL = 0
+LLC = 0
+WLC = 0
+LWC = 0
+WWC = -9.454e-17
+LWLC = 0
+WWLC = 0
+DLC = '3.70000000e-08+ddlcp_hp'
+DWC = '2.59200000e-08+ddwcp_hp'
+XPART = 0
+TOXREF = 2.35e-09
+DLCIG = 1.02e-08
+VTH0 = '-0.305+dvth0p712_hp+(mcm_PENHHP_vth0*mcmScale)'
+K1 = '0.51*dk1factorp_hp'
+K2 = '-0.1158821*dk2factorp_hp'
+K3 = 0
+K3B = 0
+W0 = 0
+DVT0 = 0
+DVT1 = 0.56
+DVT2 = 0
+DVT0W = 0
+DVT1W = 5300000
+DVT2W = 0
+DSUB = 0.56
+MINV = 0
+VOFFL = 0
+DVTP0 = 0
+DVTP1 = 0
+LPE0 = 0
+LPEB = 0
+XJ = 1.8e-08
+NGATE = 2.8e+20
+NDEP = 7.4e+17
+NSD = 1e+20
+PHIN = 0
+CDSC = 0
+CDSCB = 0
+CDSCD = 0.005035568
+CIT = 0
+VOFF = -0.1303306
+NFACTOR = 0.5046555
+ETA0 = 0.3823176
+ETAB = -0.15
+U0 = '(0.0097*du0factorp_hp)*(((1+mcm_PENHHP_u0*mcmScale)-1)+1)'
+UA = 3.4e-19
+UB = 1e-19
+UC = -7.1548571e-20
+LUC = -8.4159326e-26
+EU = 2
+VSAT = '215000*dvsatfactorp_hp'
+A0 = 0.75
+AGS = -0.1
+A1 = 0
+A2 = 0.4
+B0 = 0
+B1 = 0
+KETA = 0
+DWG = 0
+DWB = 0
+PCLM = 2.2
+PDIBLC1 = 0
+PDIBLC2 = 5.137115e-05
+PDIBLCB = -0.3660875
+DROUT = 0.56
+PVAG = 1
+DELTA = 0.01
+PSCBE1 = 2.55e+09
+PSCBE2 = 3.1e-05
+FPROUT = 0
+PDITS = 0.01
+PDITSD = 14
+PDITSL = 0
+RSH = 9
+RDSW = 511
+RSW = 256
+RDW = 256
+RDSWMIN = 0
+RDWMIN = 0
+RSWMIN = 0
+PRWG = 0.04426019
+PRWB = 0.29360737
+WR = 1
+ALPHA0 = 3.138e-09
+ALPHA1 = 0.73571
+BETA0 = 16
+AGIDL = 1.9e-06
+BGIDL = 5.357e+09
+CGIDL = 2.393
+EGIDL = -0.6972
+AIGBACC = 0.013
+BIGBACC = 0.00891
+CIGBACC = 0.0375
+NIGBACC = 10
+AIGBINV = 0.0245
+BIGBINV = 0.010197
+CIGBINV = 0
+EIGBINV = 1.1
+NIGBINV = 10
+AIGC = 0.00775
+BIGC = 0.0013
+CIGC = 2e-27
+AIGSD = 0.0062422571
+LAIGSD = -4.2079663e-10
+BIGSD = 0.0004947694
+CIGSD = 0.07079
+NIGC = 0.5
+POXEDGE = 1
+PIGCD = 1.700408
+NTOX = 1
+XRCRG1 = 12
+XRCRG2 = 1
+CGSO = '6.5e-11*dcgsofactorp_hp+dcgsop_hp'
+CGDO = '6.5e-11*dcgdofactorp_hp+dcgdop_hp'
+CGBO = 0
+CGDL = '1.4e-10*dcgdlfactorp_hp'
+CGSL = '1.4e-10*dcgslfactorp_hp'
+CLC = 0
+CLE = 0.6
+CF = '2.043195e-10*dcffactorp_hp'
+CKAPPAS = 0.6
+CKAPPAD = 0.6
+ACDE = 1
+MOIN = 15
+NOFF = 2
+VOFFCV = -0.03
+KT1 = -0.18422571
+LKT1 = 4.2079663e-08
+KT1L = 0
+KT2 = -0.04
+UTE = -1.0366143
+LUTE = -6.3119494e-07
+UA1 = 0
+UB1 = -1e-18
+UC1 = 6.8451429e-20
+LUC1 = -8.4159326e-26
+PRT = 0
+AT = 5000
+FNOIMOD = 1
+TNOIMOD = 0
+JSS = 3.36e-6
+JSWS = 1.437e-10
+JSWGS = 1.1e-8
+NJS = 1.423
+IJTHSFWD = 0.1
+JSD = 3.36e-6
+JSWD = 1.437e-10
+JSWGD = 1.1e-8
+NJD = 1.423
+IJTHDFWD = 0.1
+PBS = 0.690412
+CJS = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJS = 0.347881
+PBSWS = 0.14042
+CJSWS = '1.516703e-11*dcjfactorp_hp'
+MJSWS = 0.039289
+PBSWGS = 1.211
+CJSWGS = '293.3e-12*dcjfactorp_hp'
+MJSWGS = 900e-3
+PBD = 0.690412
+CJD = '0.0010334*dcjfactorp_hp+dcjp_hp'
+MJD = 0.347881
+PBSWD = 0.14042
+CJSWD = '1.516703e-11*dcjfactorp_hp'
+MJSWD = 0.039289
+PBSWGD = 1.211
+CJSWGD = '293.3e-12*dcjfactorp_hp'
+MJSWGD = 900e-3
+TPB = 0
+TCJ = 0
+TPBSW = 0
+TCJSW = 0
+TPBSWG = 0
+TCJSWG = 0
+XTIS = 1.5
+XTID = 1.5
+DMCG = 0
+DMCI = 0
+DMDG = 0
+DMCGT = 0
+DWJ = '2.59200000e-08+ddwjp_hp'
+XGW = 0
+XGL = 0
+RSHG = 10
+GBMIN = 1e-12
+RBPB = 50
+RBPD = 50
+RBPS = 50
+RBDB = 50
+RBSB = 50
+NGCON = 1
+XL = '0.0+dxlp_hp'
+XW = '0.0+dxwp_hp'
+LCF = '-3.66441e-18*dcffactorp_hp'
+NOIA = 2.15E+42
+NOIB = 4.0e+26
+NOIC = 8.75
+EM = 4.1e+07
+EF = 1.0
+NTNOI = 1
+LVTH0 = '0.0+dlvth0p712_hp'
+WVTH0 = '0.0+dwvth0p712_hp'
+PVTH0 = '0.0+dpvth0p712_hp'
+saref   = 1e-006          sbref   = 1e-006          wlod    = 0               kvth0   = 1e-009        
+lkvth0  = 0               wkvth0  = 0               pkvth0  = 0               llodvth = 0             
+wlodvth = 0               stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 5e-008          lku0    = 0               wku0    = 0               pku0    = 0             
+llodku0 = 0               wlodku0 = 0               kvsat   = -1              steta0  = 0             
+tku0    = 0             
+web     = 1.55e2         wec     = 2e3            kvth0we = -1.13e-2        k2we    = 3.75e-4
+ku0we   = -4.13e-3        scref   = 1e-6
+wpemod  = 1
.ENDS PENHHP_S

*** .ENDL MOS ***
