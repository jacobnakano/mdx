*simulator lang=spice

*** .LIB COMMON ***
.param
+dvth000n_hp = 0
+dvth000p_hp = 0
+du000factorn_hp = 1
+du000factorp_hp = 1
+dk100factorn_hp = 1
+dk100factorp_hp = 1
+dvth000intrn_hp = 2.27m
+dvth000intrp_hp = 2.40m

*** .ENDL COMMON ***

