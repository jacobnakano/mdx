*simulator lang=spice
*** .LIB COMMON_DVTH ***
.param
+dvth0n001_hp = '1.7123e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n001_hp = '8.4413e-09*dvth0intrn_hp'
+dwvth0n001_hp = '5.3948e-06*dvth0intrn_hp'
+dpvth0n001_hp = '2.6595e-13*dvth0intrn_hp'
+dvth0n101_hp = '4.6309e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n101_hp = '2.2829e-08*dvth0intrn_hp'
+dwvth0n101_hp = '2.4972e-06*dvth0intrn_hp'
+dpvth0n101_hp = '1.2311e-13*dvth0intrn_hp'
+dvth0n201_hp = '8.4150e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n201_hp = '4.1484e-08*dvth0intrn_hp'
+dwvth0n201_hp = '1.3889e-06*dvth0intrn_hp'
+dpvth0n201_hp = '6.8467e-14*dvth0intrn_hp'
+dvth0n301_hp = '1.3885e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n301_hp = '6.8451e-08*dvth0intrn_hp'
+dwvth0n301_hp = '8.8012e-07*dvth0intrn_hp'
+dpvth0n301_hp = '4.3387e-14*dvth0intrn_hp'
+dvth0n401_hp = '2.0865e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n401_hp = '1.0286e-07*dvth0intrn_hp'
+dwvth0n401_hp = '5.7859e-07*dvth0intrn_hp'
+dpvth0n401_hp = '2.8523e-14*dvth0intrn_hp'
+dvth0n501_hp = '3.0840e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n501_hp = '1.5203e-07*dvth0intrn_hp'
+dwvth0n501_hp = '4.0104e-07*dvth0intrn_hp'
+dpvth0n501_hp = '1.9770e-14*dvth0intrn_hp'
+dvth0n601_hp = '3.9311e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n601_hp = '1.9379e-07*dvth0intrn_hp'
+dwvth0n601_hp = '3.2057e-07*dvth0intrn_hp'
+dpvth0n601_hp = '1.5803e-14*dvth0intrn_hp'
+dvth0n002_hp = '1.6704e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n002_hp = '8.6544e-09*dvth0intrn_hp'
+dwvth0n002_hp = '5.2627e-06*dvth0intrn_hp'
+dpvth0n002_hp = '2.7266e-13*dvth0intrn_hp'
+dvth0n102_hp = '4.5175e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n102_hp = '2.3405e-08*dvth0intrn_hp'
+dwvth0n102_hp = '2.4361e-06*dvth0intrn_hp'
+dpvth0n102_hp = '1.2621e-13*dvth0intrn_hp'
+dvth0n202_hp = '8.2090e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n202_hp = '4.2531e-08*dvth0intrn_hp'
+dwvth0n202_hp = '1.3548e-06*dvth0intrn_hp'
+dpvth0n202_hp = '7.0195e-14*dvth0intrn_hp'
+dvth0n302_hp = '1.3545e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n302_hp = '7.0179e-08*dvth0intrn_hp'
+dwvth0n302_hp = '8.5856e-07*dvth0intrn_hp'
+dpvth0n302_hp = '4.4482e-14*dvth0intrn_hp'
+dvth0n402_hp = '2.0354e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n402_hp = '1.0546e-07*dvth0intrn_hp'
+dwvth0n402_hp = '5.6442e-07*dvth0intrn_hp'
+dpvth0n402_hp = '2.9243e-14*dvth0intrn_hp'
+dvth0n502_hp = '3.0085e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n502_hp = '1.5587e-07*dvth0intrn_hp'
+dwvth0n502_hp = '3.9122e-07*dvth0intrn_hp'
+dpvth0n502_hp = '2.0269e-14*dvth0intrn_hp'
+dvth0n602_hp = '3.8348e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n602_hp = '1.9868e-07*dvth0intrn_hp'
+dwvth0n602_hp = '3.1272e-07*dvth0intrn_hp'
+dpvth0n602_hp = '1.6202e-14*dvth0intrn_hp'
+dvth0n003_hp = '1.6099e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n003_hp = '8.9737e-09*dvth0intrn_hp'
+dwvth0n003_hp = '5.0722e-06*dvth0intrn_hp'
+dpvth0n003_hp = '2.8272e-13*dvth0intrn_hp'
+dvth0n103_hp = '4.3540e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n103_hp = '2.4269e-08*dvth0intrn_hp'
+dwvth0n103_hp = '2.3479e-06*dvth0intrn_hp'
+dpvth0n103_hp = '1.3087e-13*dvth0intrn_hp'
+dvth0n203_hp = '7.9119e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n203_hp = '4.4100e-08*dvth0intrn_hp'
+dwvth0n203_hp = '1.3058e-06*dvth0intrn_hp'
+dpvth0n203_hp = '7.2785e-14*dvth0intrn_hp'
+dvth0n303_hp = '1.3055e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n303_hp = '7.2768e-08*dvth0intrn_hp'
+dwvth0n303_hp = '8.2749e-07*dvth0intrn_hp'
+dpvth0n303_hp = '4.6124e-14*dvth0intrn_hp'
+dvth0n403_hp = '1.9617e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n403_hp = '1.0935e-07*dvth0intrn_hp'
+dwvth0n403_hp = '5.4400e-07*dvth0intrn_hp'
+dpvth0n403_hp = '3.0322e-14*dvth0intrn_hp'
+dvth0n503_hp = '2.8996e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n503_hp = '1.6162e-07*dvth0intrn_hp'
+dwvth0n503_hp = '3.7706e-07*dvth0intrn_hp'
+dpvth0n503_hp = '2.1017e-14*dvth0intrn_hp'
+dvth0n603_hp = '3.6960e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n603_hp = '2.0601e-07*dvth0intrn_hp'
+dwvth0n603_hp = '3.0140e-07*dvth0intrn_hp'
+dpvth0n603_hp = '1.6800e-14*dvth0intrn_hp'
+dvth0n004_hp = '1.5612e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n004_hp = '9.2606e-09*dvth0intrn_hp'
+dwvth0n004_hp = '4.9186e-06*dvth0intrn_hp'
+dpvth0n004_hp = '2.9176e-13*dvth0intrn_hp'
+dvth0n104_hp = '4.2221e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n104_hp = '2.5045e-08*dvth0intrn_hp'
+dwvth0n104_hp = '2.2768e-06*dvth0intrn_hp'
+dpvth0n104_hp = '1.3505e-13*dvth0intrn_hp'
+dvth0n204_hp = '7.6722e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n204_hp = '4.5510e-08*dvth0intrn_hp'
+dwvth0n204_hp = '1.2663e-06*dvth0intrn_hp'
+dpvth0n204_hp = '7.5112e-14*dvth0intrn_hp'
+dvth0n304_hp = '1.2660e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n304_hp = '7.5094e-08*dvth0intrn_hp'
+dwvth0n304_hp = '8.0242e-07*dvth0intrn_hp'
+dpvth0n304_hp = '4.7598e-14*dvth0intrn_hp'
+dvth0n404_hp = '1.9023e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n404_hp = '1.1284e-07*dvth0intrn_hp'
+dwvth0n404_hp = '5.2752e-07*dvth0intrn_hp'
+dpvth0n404_hp = '3.1291e-14*dvth0intrn_hp'
+dvth0n504_hp = '2.8118e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n504_hp = '1.6679e-07*dvth0intrn_hp'
+dwvth0n504_hp = '3.6564e-07*dvth0intrn_hp'
+dpvth0n504_hp = '2.1689e-14*dvth0intrn_hp'
+dvth0n604_hp = '3.5840e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n604_hp = '2.1260e-07*dvth0intrn_hp'
+dwvth0n604_hp = '2.9227e-07*dvth0intrn_hp'
+dpvth0n604_hp = '1.7337e-14*dvth0intrn_hp'
+dvth0n005_hp = '1.5175e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n005_hp = '9.5219e-09*dvth0intrn_hp'
+dwvth0n005_hp = '4.7809e-06*dvth0intrn_hp'
+dpvth0n005_hp = '2.9999e-13*dvth0intrn_hp'
+dvth0n105_hp = '4.1040e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n105_hp = '2.5752e-08*dvth0intrn_hp'
+dwvth0n105_hp = '2.2131e-06*dvth0intrn_hp'
+dpvth0n105_hp = '1.3887e-13*dvth0intrn_hp'
+dvth0n205_hp = '7.4575e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n205_hp = '4.6794e-08*dvth0intrn_hp'
+dwvth0n205_hp = '1.2308e-06*dvth0intrn_hp'
+dpvth0n205_hp = '7.7232e-14*dvth0intrn_hp'
+dvth0n305_hp = '1.2305e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n305_hp = '7.7214e-08*dvth0intrn_hp'
+dwvth0n305_hp = '7.7997e-07*dvth0intrn_hp'
+dpvth0n305_hp = '4.8942e-14*dvth0intrn_hp'
+dvth0n405_hp = '1.8491e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n405_hp = '1.1603e-07*dvth0intrn_hp'
+dwvth0n405_hp = '5.1275e-07*dvth0intrn_hp'
+dpvth0n405_hp = '3.2174e-14*dvth0intrn_hp'
+dvth0n505_hp = '2.7331e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n505_hp = '1.7150e-07*dvth0intrn_hp'
+dwvth0n505_hp = '3.5540e-07*dvth0intrn_hp'
+dpvth0n505_hp = '2.2301e-14*dvth0intrn_hp'
+dvth0n605_hp = '3.4837e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n605_hp = '2.1860e-07*dvth0intrn_hp'
+dwvth0n605_hp = '2.8409e-07*dvth0intrn_hp'
+dpvth0n605_hp = '1.7826e-14*dvth0intrn_hp'
+dvth0n006_hp = '1.4602e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n006_hp = '9.8989e-09*dvth0intrn_hp'
+dwvth0n006_hp = '4.6005e-06*dvth0intrn_hp'
+dpvth0n006_hp = '3.1187e-13*dvth0intrn_hp'
+dvth0n106_hp = '3.9491e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n106_hp = '2.6771e-08*dvth0intrn_hp'
+dwvth0n106_hp = '2.1295e-06*dvth0intrn_hp'
+dpvth0n106_hp = '1.4436e-13*dvth0intrn_hp'
+dvth0n206_hp = '7.1760e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n206_hp = '4.8647e-08*dvth0intrn_hp'
+dwvth0n206_hp = '1.1844e-06*dvth0intrn_hp'
+dpvth0n206_hp = '8.0289e-14*dvth0intrn_hp'
+dvth0n306_hp = '1.1841e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n306_hp = '8.0270e-08*dvth0intrn_hp'
+dwvth0n306_hp = '7.5053e-07*dvth0intrn_hp'
+dpvth0n306_hp = '5.0879e-14*dvth0intrn_hp'
+dvth0n406_hp = '1.7793e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n406_hp = '1.2062e-07*dvth0intrn_hp'
+dwvth0n406_hp = '4.9340e-07*dvth0intrn_hp'
+dpvth0n406_hp = '3.3448e-14*dvth0intrn_hp'
+dvth0n506_hp = '2.6299e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n506_hp = '1.7828e-07*dvth0intrn_hp'
+dwvth0n506_hp = '3.4199e-07*dvth0intrn_hp'
+dpvth0n506_hp = '2.3184e-14*dvth0intrn_hp'
+dvth0n606_hp = '3.3523e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n606_hp = '2.2725e-07*dvth0intrn_hp'
+dwvth0n606_hp = '2.7337e-07*dvth0intrn_hp'
+dpvth0n606_hp = '1.8532e-14*dvth0intrn_hp'
+dvth0n007_hp = '1.4204e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n007_hp = '1.0177e-08*dvth0intrn_hp'
+dwvth0n007_hp = '4.4751e-06*dvth0intrn_hp'
+dpvth0n007_hp = '3.2062e-13*dvth0intrn_hp'
+dvth0n107_hp = '3.8415e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n107_hp = '2.7523e-08*dvth0intrn_hp'
+dwvth0n107_hp = '2.0715e-06*dvth0intrn_hp'
+dpvth0n107_hp = '1.4842e-13*dvth0intrn_hp'
+dvth0n207_hp = '6.9805e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n207_hp = '5.0012e-08*dvth0intrn_hp'
+dwvth0n207_hp = '1.1521e-06*dvth0intrn_hp'
+dpvth0n207_hp = '8.2543e-14*dvth0intrn_hp'
+dvth0n307_hp = '1.1518e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n307_hp = '8.2524e-08*dvth0intrn_hp'
+dwvth0n307_hp = '7.3008e-07*dvth0intrn_hp'
+dpvth0n307_hp = '5.2307e-14*dvth0intrn_hp'
+dvth0n407_hp = '1.7308e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n407_hp = '1.2401e-07*dvth0intrn_hp'
+dwvth0n407_hp = '4.7995e-07*dvth0intrn_hp'
+dpvth0n407_hp = '3.4387e-14*dvth0intrn_hp'
+dvth0n507_hp = '2.5582e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n507_hp = '1.8329e-07*dvth0intrn_hp'
+dwvth0n507_hp = '3.3267e-07*dvth0intrn_hp'
+dpvth0n507_hp = '2.3835e-14*dvth0intrn_hp'
+dvth0n607_hp = '3.2609e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n607_hp = '2.3363e-07*dvth0intrn_hp'
+dwvth0n607_hp = '2.6592e-07*dvth0intrn_hp'
+dpvth0n607_hp = '1.9052e-14*dvth0intrn_hp'
+dvth0n008_hp = '1.3441e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n008_hp = '1.0738e-08*dvth0intrn_hp'
+dwvth0n008_hp = '4.2345e-06*dvth0intrn_hp'
+dpvth0n008_hp = '3.3831e-13*dvth0intrn_hp'
+dvth0n108_hp = '3.6349e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n108_hp = '2.9041e-08*dvth0intrn_hp'
+dwvth0n108_hp = '1.9601e-06*dvth0intrn_hp'
+dpvth0n108_hp = '1.5660e-13*dvth0intrn_hp'
+dvth0n208_hp = '6.6052e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n208_hp = '5.2771e-08*dvth0intrn_hp'
+dwvth0n208_hp = '1.0902e-06*dvth0intrn_hp'
+dpvth0n208_hp = '8.7096e-14*dvth0intrn_hp'
+dvth0n308_hp = '1.0899e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n308_hp = '8.7076e-08*dvth0intrn_hp'
+dwvth0n308_hp = '6.9083e-07*dvth0intrn_hp'
+dpvth0n308_hp = '5.5193e-14*dvth0intrn_hp'
+dvth0n408_hp = '1.6378e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n408_hp = '1.3085e-07*dvth0intrn_hp'
+dwvth0n408_hp = '4.5415e-07*dvth0intrn_hp'
+dpvth0n408_hp = '3.6284e-14*dvth0intrn_hp'
+dvth0n508_hp = '2.4207e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n508_hp = '1.9340e-07*dvth0intrn_hp'
+dwvth0n508_hp = '3.1479e-07*dvth0intrn_hp'
+dpvth0n508_hp = '2.5149e-14*dvth0intrn_hp'
+dvth0n608_hp = '3.0856e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n608_hp = '2.4652e-07*dvth0intrn_hp'
+dwvth0n608_hp = '2.5162e-07*dvth0intrn_hp'
+dpvth0n608_hp = '2.0103e-14*dvth0intrn_hp'
+dvth0n009_hp = '1.2759e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n009_hp = '1.1330e-08*dvth0intrn_hp'
+dwvth0n009_hp = '4.0198e-06*dvth0intrn_hp'
+dpvth0n009_hp = '3.5695e-13*dvth0intrn_hp'
+dvth0n109_hp = '3.4506e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n109_hp = '3.0641e-08*dvth0intrn_hp'
+dwvth0n109_hp = '1.8608e-06*dvth0intrn_hp'
+dpvth0n109_hp = '1.6523e-13*dvth0intrn_hp'
+dvth0n209_hp = '6.2703e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n209_hp = '5.5679e-08*dvth0intrn_hp'
+dwvth0n209_hp = '1.0349e-06*dvth0intrn_hp'
+dpvth0n209_hp = '9.1895e-14*dvth0intrn_hp'
+dvth0n309_hp = '1.0346e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n309_hp = '9.1874e-08*dvth0intrn_hp'
+dwvth0n309_hp = '6.5580e-07*dvth0intrn_hp'
+dpvth0n309_hp = '5.8234e-14*dvth0intrn_hp'
+dvth0n409_hp = '1.5547e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n409_hp = '1.3806e-07*dvth0intrn_hp'
+dwvth0n409_hp = '4.3113e-07*dvth0intrn_hp'
+dpvth0n409_hp = '3.8283e-14*dvth0intrn_hp'
+dvth0n509_hp = '2.2980e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n509_hp = '2.0406e-07*dvth0intrn_hp'
+dwvth0n509_hp = '2.9883e-07*dvth0intrn_hp'
+dpvth0n509_hp = '2.6535e-14*dvth0intrn_hp'
+dvth0n609_hp = '2.9292e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n609_hp = '2.6010e-07*dvth0intrn_hp'
+dwvth0n609_hp = '2.3887e-07*dvth0intrn_hp'
+dpvth0n609_hp = '2.1211e-14*dvth0intrn_hp'
+dvth0n010_hp = '1.2481e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n010_hp = '1.1582e-08*dvth0intrn_hp'
+dwvth0n010_hp = '3.9322e-06*dvth0intrn_hp'
+dpvth0n010_hp = '3.6491e-13*dvth0intrn_hp'
+dvth0n110_hp = '3.3755e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n110_hp = '3.1324e-08*dvth0intrn_hp'
+dwvth0n110_hp = '1.8202e-06*dvth0intrn_hp'
+dpvth0n110_hp = '1.6891e-13*dvth0intrn_hp'
+dvth0n210_hp = '6.1337e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n210_hp = '5.6920e-08*dvth0intrn_hp'
+dwvth0n210_hp = '1.0123e-06*dvth0intrn_hp'
+dpvth0n210_hp = '9.3943e-14*dvth0intrn_hp'
+dvth0n310_hp = '1.0121e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n310_hp = '9.3921e-08*dvth0intrn_hp'
+dwvth0n310_hp = '6.4151e-07*dvth0intrn_hp'
+dpvth0n310_hp = '5.9531e-14*dvth0intrn_hp'
+dvth0n410_hp = '1.5208e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n410_hp = '1.4113e-07*dvth0intrn_hp'
+dwvth0n410_hp = '4.2173e-07*dvth0intrn_hp'
+dpvth0n410_hp = '3.9136e-14*dvth0intrn_hp'
+dvth0n510_hp = '2.2479e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n510_hp = '2.0860e-07*dvth0intrn_hp'
+dwvth0n510_hp = '2.9232e-07*dvth0intrn_hp'
+dpvth0n510_hp = '2.7126e-14*dvth0intrn_hp'
+dvth0n610_hp = '2.8653e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n610_hp = '2.6590e-07*dvth0intrn_hp'
+dwvth0n610_hp = '2.3366e-07*dvth0intrn_hp'
+dpvth0n610_hp = '2.1683e-14*dvth0intrn_hp'
+dvth0n011_hp = '1.0862e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n011_hp = '1.3118e-08*dvth0intrn_hp'
+dwvth0n011_hp = '3.4221e-06*dvth0intrn_hp'
+dpvth0n011_hp = '4.1328e-13*dvth0intrn_hp'
+dvth0n111_hp = '2.9375e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n111_hp = '3.5476e-08*dvth0intrn_hp'
+dwvth0n111_hp = '1.5841e-06*dvth0intrn_hp'
+dpvth0n111_hp = '1.9131e-13*dvth0intrn_hp'
+dvth0n211_hp = '5.3379e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n211_hp = '6.4465e-08*dvth0intrn_hp'
+dwvth0n211_hp = '8.8099e-07*dvth0intrn_hp'
+dpvth0n211_hp = '1.0640e-13*dvth0intrn_hp'
+dvth0n311_hp = '8.8079e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n311_hp = '1.0637e-07*dvth0intrn_hp'
+dwvth0n311_hp = '5.5828e-07*dvth0intrn_hp'
+dpvth0n311_hp = '6.7423e-14*dvth0intrn_hp'
+dvth0n411_hp = '1.3235e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n411_hp = '1.5984e-07*dvth0intrn_hp'
+dwvth0n411_hp = '3.6702e-07*dvth0intrn_hp'
+dpvth0n411_hp = '4.4324e-14*dvth0intrn_hp'
+dvth0n511_hp = '1.9563e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n511_hp = '2.3626e-07*dvth0intrn_hp'
+dwvth0n511_hp = '2.5439e-07*dvth0intrn_hp'
+dpvth0n511_hp = '3.0722e-14*dvth0intrn_hp'
+dvth0n611_hp = '2.4936e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n611_hp = '3.0115e-07*dvth0intrn_hp'
+dwvth0n611_hp = '2.0335e-07*dvth0intrn_hp'
+dpvth0n611_hp = '2.4558e-14*dvth0intrn_hp'
+dvth0n012_hp = '9.6327e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n012_hp = '1.5008e-08*dvth0intrn_hp'
+dwvth0n012_hp = '3.0348e-06*dvth0intrn_hp'
+dpvth0n012_hp = '4.7285e-13*dvth0intrn_hp'
+dvth0n112_hp = '2.6051e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n112_hp = '4.0589e-08*dvth0intrn_hp'
+dwvth0n112_hp = '1.4048e-06*dvth0intrn_hp'
+dpvth0n112_hp = '2.1888e-13*dvth0intrn_hp'
+dvth0n212_hp = '4.7338e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n212_hp = '7.3757e-08*dvth0intrn_hp'
+dwvth0n212_hp = '7.8130e-07*dvth0intrn_hp'
+dpvth0n212_hp = '1.2173e-13*dvth0intrn_hp'
+dvth0n312_hp = '7.8112e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n312_hp = '1.2170e-07*dvth0intrn_hp'
+dwvth0n312_hp = '4.9511e-07*dvth0intrn_hp'
+dpvth0n312_hp = '7.7141e-14*dvth0intrn_hp'
+dvth0n412_hp = '1.1738e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n412_hp = '1.8288e-07*dvth0intrn_hp'
+dwvth0n412_hp = '3.2548e-07*dvth0intrn_hp'
+dpvth0n412_hp = '5.0713e-14*dvth0intrn_hp'
+dvth0n512_hp = '1.7349e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n512_hp = '2.7031e-07*dvth0intrn_hp'
+dwvth0n512_hp = '2.2560e-07*dvth0intrn_hp'
+dpvth0n512_hp = '3.5151e-14*dvth0intrn_hp'
+dvth0n612_hp = '2.2114e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n612_hp = '3.4455e-07*dvth0intrn_hp'
+dwvth0n612_hp = '1.8033e-07*dvth0intrn_hp'
+dpvth0n612_hp = '2.8097e-14*dvth0intrn_hp'
+dvth0n013_hp = '9.5113e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n013_hp = '1.5200e-08*dvth0intrn_hp'
+dwvth0n013_hp = '2.9966e-06*dvth0intrn_hp'
+dpvth0n013_hp = '4.7888e-13*dvth0intrn_hp'
+dvth0n113_hp = '2.5723e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n113_hp = '4.1107e-08*dvth0intrn_hp'
+dwvth0n113_hp = '1.3871e-06*dvth0intrn_hp'
+dpvth0n113_hp = '2.2167e-13*dvth0intrn_hp'
+dvth0n213_hp = '4.6742e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n213_hp = '7.4698e-08*dvth0intrn_hp'
+dwvth0n213_hp = '7.7146e-07*dvth0intrn_hp'
+dpvth0n213_hp = '1.2328e-13*dvth0intrn_hp'
+dvth0n313_hp = '7.7128e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n313_hp = '1.2326e-07*dvth0intrn_hp'
+dwvth0n313_hp = '4.8887e-07*dvth0intrn_hp'
+dpvth0n313_hp = '7.8125e-14*dvth0intrn_hp'
+dvth0n413_hp = '1.1590e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n413_hp = '1.8521e-07*dvth0intrn_hp'
+dwvth0n413_hp = '3.2139e-07*dvth0intrn_hp'
+dpvth0n413_hp = '5.1360e-14*dvth0intrn_hp'
+dvth0n513_hp = '1.7130e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n513_hp = '2.7376e-07*dvth0intrn_hp'
+dwvth0n513_hp = '2.2276e-07*dvth0intrn_hp'
+dpvth0n513_hp = '3.5599e-14*dvth0intrn_hp'
+dvth0n613_hp = '2.1835e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n613_hp = '3.4895e-07*dvth0intrn_hp'
+dwvth0n613_hp = '1.7806e-07*dvth0intrn_hp'
+dpvth0n613_hp = '2.8456e-14*dvth0intrn_hp'
+dvth0n014_hp = '8.4394e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n014_hp = '1.6934e-08*dvth0intrn_hp'
+dwvth0n014_hp = '2.6589e-06*dvth0intrn_hp'
+dpvth0n014_hp = '5.3353e-13*dvth0intrn_hp'
+dvth0n114_hp = '2.2824e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n114_hp = '4.5798e-08*dvth0intrn_hp'
+dwvth0n114_hp = '1.2308e-06*dvth0intrn_hp'
+dpvth0n114_hp = '2.4697e-13*dvth0intrn_hp'
+dvth0n214_hp = '4.1474e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n214_hp = '8.3222e-08*dvth0intrn_hp'
+dwvth0n214_hp = '6.8451e-07*dvth0intrn_hp'
+dpvth0n214_hp = '1.3735e-13*dvth0intrn_hp'
+dvth0n314_hp = '6.8435e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n314_hp = '1.3732e-07*dvth0intrn_hp'
+dwvth0n314_hp = '4.3377e-07*dvth0intrn_hp'
+dpvth0n314_hp = '8.7041e-14*dvth0intrn_hp'
+dvth0n414_hp = '1.0284e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n414_hp = '2.0635e-07*dvth0intrn_hp'
+dwvth0n414_hp = '2.8516e-07*dvth0intrn_hp'
+dpvth0n414_hp = '5.7221e-14*dvth0intrn_hp'
+dvth0n514_hp = '1.5200e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n514_hp = '3.0500e-07*dvth0intrn_hp'
+dwvth0n514_hp = '1.9766e-07*dvth0intrn_hp'
+dpvth0n514_hp = '3.9661e-14*dvth0intrn_hp'
+dvth0n614_hp = '1.9375e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n614_hp = '3.8877e-07*dvth0intrn_hp'
+dwvth0n614_hp = '1.5800e-07*dvth0intrn_hp'
+dpvth0n614_hp = '3.1703e-14*dvth0intrn_hp'
+dvth0n015_hp = '7.5923e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n015_hp = '1.9042e-08*dvth0intrn_hp'
+dwvth0n015_hp = '2.3920e-06*dvth0intrn_hp'
+dpvth0n015_hp = '5.9994e-13*dvth0intrn_hp'
+dvth0n115_hp = '2.0533e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n115_hp = '5.1499e-08*dvth0intrn_hp'
+dwvth0n115_hp = '1.1072e-06*dvth0intrn_hp'
+dpvth0n115_hp = '2.7771e-13*dvth0intrn_hp'
+dvth0n215_hp = '3.7311e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n215_hp = '9.3581e-08*dvth0intrn_hp'
+dwvth0n215_hp = '6.1580e-07*dvth0intrn_hp'
+dpvth0n215_hp = '1.5445e-13*dvth0intrn_hp'
+dvth0n315_hp = '6.1566e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n315_hp = '1.5441e-07*dvth0intrn_hp'
+dwvth0n315_hp = '3.9023e-07*dvth0intrn_hp'
+dpvth0n315_hp = '9.7875e-14*dvth0intrn_hp'
+dvth0n415_hp = '9.2513e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n415_hp = '2.3203e-07*dvth0intrn_hp'
+dwvth0n415_hp = '2.5654e-07*dvth0intrn_hp'
+dpvth0n415_hp = '6.4343e-14*dvth0intrn_hp'
+dvth0n515_hp = '1.3674e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n515_hp = '3.4296e-07*dvth0intrn_hp'
+dwvth0n515_hp = '1.7782e-07*dvth0intrn_hp'
+dpvth0n515_hp = '4.4598e-14*dvth0intrn_hp'
+dvth0n615_hp = '1.7430e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n615_hp = '4.3716e-07*dvth0intrn_hp'
+dwvth0n615_hp = '1.4214e-07*dvth0intrn_hp'
+dpvth0n615_hp = '3.5649e-14*dvth0intrn_hp'
+dvth0n016_hp = '7.5324e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n016_hp = '1.9194e-08*dvth0intrn_hp'
+dwvth0n016_hp = '2.3731e-06*dvth0intrn_hp'
+dpvth0n016_hp = '6.0470e-13*dvth0intrn_hp'
+dvth0n116_hp = '2.0371e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n116_hp = '5.1908e-08*dvth0intrn_hp'
+dwvth0n116_hp = '1.0985e-06*dvth0intrn_hp'
+dpvth0n116_hp = '2.7991e-13*dvth0intrn_hp'
+dvth0n216_hp = '3.7017e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n216_hp = '9.4324e-08*dvth0intrn_hp'
+dwvth0n216_hp = '6.1095e-07*dvth0intrn_hp'
+dpvth0n216_hp = '1.5568e-13*dvth0intrn_hp'
+dvth0n316_hp = '6.1081e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n316_hp = '1.5564e-07*dvth0intrn_hp'
+dwvth0n316_hp = '3.8716e-07*dvth0intrn_hp'
+dpvth0n316_hp = '9.8652e-14*dvth0intrn_hp'
+dvth0n416_hp = '9.1784e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n416_hp = '2.3388e-07*dvth0intrn_hp'
+dwvth0n416_hp = '2.5452e-07*dvth0intrn_hp'
+dpvth0n416_hp = '6.4854e-14*dvth0intrn_hp'
+dvth0n516_hp = '1.3566e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n516_hp = '3.4569e-07*dvth0intrn_hp'
+dwvth0n516_hp = '1.7641e-07*dvth0intrn_hp'
+dpvth0n516_hp = '4.4952e-14*dvth0intrn_hp'
+dvth0n616_hp = '1.7292e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n616_hp = '4.4063e-07*dvth0intrn_hp'
+dwvth0n616_hp = '1.4102e-07*dvth0intrn_hp'
+dpvth0n616_hp = '3.5933e-14*dvth0intrn_hp'
+dvth0n017_hp = '5.1194e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n017_hp = '2.5391e-08*dvth0intrn_hp'
+dwvth0n017_hp = '1.6129e-06*dvth0intrn_hp'
+dpvth0n017_hp = '7.9995e-13*dvth0intrn_hp'
+dvth0n117_hp = '1.3845e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n117_hp = '6.8668e-08*dvth0intrn_hp'
+dwvth0n117_hp = '7.4660e-07*dvth0intrn_hp'
+dpvth0n117_hp = '3.7029e-13*dvth0intrn_hp'
+dvth0n217_hp = '2.5159e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n217_hp = '1.2478e-07*dvth0intrn_hp'
+dwvth0n217_hp = '4.1523e-07*dvth0intrn_hp'
+dpvth0n217_hp = '2.0594e-13*dvth0intrn_hp'
+dvth0n317_hp = '4.1513e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n317_hp = '2.0589e-07*dvth0intrn_hp'
+dwvth0n317_hp = '2.6313e-07*dvth0intrn_hp'
+dpvth0n317_hp = '1.3051e-13*dvth0intrn_hp'
+dvth0n417_hp = '6.2381e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n417_hp = '3.0939e-07*dvth0intrn_hp'
+dwvth0n417_hp = '1.7298e-07*dvth0intrn_hp'
+dpvth0n417_hp = '8.5794e-14*dvth0intrn_hp'
+dvth0n517_hp = '9.2203e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n517_hp = '4.5730e-07*dvth0intrn_hp'
+dwvth0n517_hp = '1.1990e-07*dvth0intrn_hp'
+dpvth0n517_hp = '5.9467e-14*dvth0intrn_hp'
+dvth0n617_hp = '1.1753e+00*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n617_hp = '5.8290e-07*dvth0intrn_hp'
+dwvth0n617_hp = '9.5841e-08*dvth0intrn_hp'
+dpvth0n617_hp = '4.7534e-14*dvth0intrn_hp'
+dvth0n018_hp = '2.8181e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n018_hp = '4.7433e-08*dvth0intrn_hp'
+dwvth0n018_hp = '8.8785e-07*dvth0intrn_hp'
+dpvth0n018_hp = '1.4944e-12*dvth0intrn_hp'
+dvth0n118_hp = '7.6214e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n118_hp = '1.2828e-07*dvth0intrn_hp'
+dwvth0n118_hp = '4.1098e-07*dvth0intrn_hp'
+dpvth0n118_hp = '6.9175e-13*dvth0intrn_hp'
+dvth0n218_hp = '1.3849e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n218_hp = '2.3310e-07*dvth0intrn_hp'
+dwvth0n218_hp = '2.2857e-07*dvth0intrn_hp'
+dpvth0n218_hp = '3.8473e-13*dvth0intrn_hp'
+dvth0n318_hp = '2.2852e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n318_hp = '3.8464e-07*dvth0intrn_hp'
+dwvth0n318_hp = '1.4485e-07*dvth0intrn_hp'
+dpvth0n318_hp = '2.4380e-13*dvth0intrn_hp'
+dvth0n418_hp = '3.4339e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n418_hp = '5.7798e-07*dvth0intrn_hp'
+dwvth0n418_hp = '9.5222e-08*dvth0intrn_hp'
+dpvth0n418_hp = '1.6028e-13*dvth0intrn_hp'
+dvth0n518_hp = '5.0755e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n518_hp = '8.5430e-07*dvth0intrn_hp'
+dwvth0n518_hp = '6.6001e-08*dvth0intrn_hp'
+dpvth0n518_hp = '1.1109e-13*dvth0intrn_hp'
+dvth0n618_hp = '6.4696e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n618_hp = '1.0889e-06*dvth0intrn_hp'
+dwvth0n618_hp = '5.2758e-08*dvth0intrn_hp'
+dpvth0n618_hp = '8.8800e-14*dvth0intrn_hp'
+dvth0n019_hp = '1.5598e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n019_hp = '8.4651e-08*dvth0intrn_hp'
+dwvth0n019_hp = '4.9142e-07*dvth0intrn_hp'
+dpvth0n019_hp = '2.6670e-12*dvth0intrn_hp'
+dvth0n119_hp = '4.2184e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n119_hp = '2.2894e-07*dvth0intrn_hp'
+dwvth0n119_hp = '2.2748e-07*dvth0intrn_hp'
+dpvth0n119_hp = '1.2345e-12*dvth0intrn_hp'
+dvth0n219_hp = '7.6654e-02*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n219_hp = '4.1601e-07*dvth0intrn_hp'
+dwvth0n219_hp = '1.2651e-07*dvth0intrn_hp'
+dpvth0n219_hp = '6.8660e-13*dvth0intrn_hp'
+dvth0n319_hp = '1.2648e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n319_hp = '6.8644e-07*dvth0intrn_hp'
+dwvth0n319_hp = '8.0171e-08*dvth0intrn_hp'
+dpvth0n319_hp = '4.3510e-13*dvth0intrn_hp'
+dvth0n419_hp = '1.9006e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n419_hp = '1.0315e-06*dvth0intrn_hp'
+dwvth0n419_hp = '5.2705e-08*dvth0intrn_hp'
+dpvth0n419_hp = '2.8603e-13*dvth0intrn_hp'
+dvth0n519_hp = '2.8093e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n519_hp = '1.5246e-06*dvth0intrn_hp'
+dwvth0n519_hp = '3.6531e-08*dvth0intrn_hp'
+dpvth0n519_hp = '1.9826e-13*dvth0intrn_hp'
+dvth0n619_hp = '3.5809e-01*dvth0intrn_hp+dvth0shiftn_hp'
+dlvth0n619_hp = '1.9434e-06*dvth0intrn_hp'
+dwvth0n619_hp = '2.9201e-08*dvth0intrn_hp'
+dpvth0n619_hp = '1.5848e-13*dvth0intrn_hp'
+dvth0p001_hp = '1.6798e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p001_hp = '8.5938e-09*dvth0intrp_hp'
+dwvth0p001_hp = '5.3047e-06*dvth0intrp_hp'
+dpvth0p001_hp = '2.7138e-13*dvth0intrp_hp'
+dvth0p101_hp = '4.5284e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p101_hp = '2.3167e-08*dvth0intrp_hp'
+dwvth0p101_hp = '2.4646e-06*dvth0intrp_hp'
+dpvth0p101_hp = '1.2609e-13*dvth0intrp_hp'
+dvth0p201_hp = '8.1579e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p201_hp = '4.1735e-08*dvth0intrp_hp'
+dwvth0p201_hp = '1.3863e-06*dvth0intrp_hp'
+dpvth0p201_hp = '7.0922e-14*dvth0intrp_hp'
+dvth0p301_hp = '1.3201e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p301_hp = '6.7537e-08*dvth0intrp_hp'
+dwvth0p301_hp = '8.9607e-07*dvth0intrp_hp'
+dpvth0p301_hp = '4.5842e-14*dvth0intrp_hp'
+dvth0p401_hp = '1.9096e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p401_hp = '9.7694e-08*dvth0intrp_hp'
+dwvth0p401_hp = '6.1666e-07*dvth0intrp_hp'
+dpvth0p401_hp = '3.1548e-14*dvth0intrp_hp'
+dvth0p501_hp = '2.6340e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p501_hp = '1.3475e-07*dvth0intrp_hp'
+dwvth0p501_hp = '4.5729e-07*dvth0intrp_hp'
+dpvth0p501_hp = '2.3395e-14*dvth0intrp_hp'
+dvth0p601_hp = '3.1362e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p601_hp = '1.6045e-07*dvth0intrp_hp'
+dwvth0p601_hp = '3.8849e-07*dvth0intrp_hp'
+dpvth0p601_hp = '1.9875e-14*dvth0intrp_hp'
+dvth0p701_hp = '3.3796e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p701_hp = '1.7290e-07*dvth0intrp_hp'
+dwvth0p701_hp = '3.6123e-07*dvth0intrp_hp'
+dpvth0p701_hp = '1.8480e-14*dvth0intrp_hp'
+dvth0p002_hp = '1.6125e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p002_hp = '8.9471e-09*dvth0intrp_hp'
+dwvth0p002_hp = '5.0920e-06*dvth0intrp_hp'
+dpvth0p002_hp = '2.8254e-13*dvth0intrp_hp'
+dvth0p102_hp = '4.3469e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p102_hp = '2.4119e-08*dvth0intrp_hp'
+dwvth0p102_hp = '2.3658e-06*dvth0intrp_hp'
+dpvth0p102_hp = '1.3127e-13*dvth0intrp_hp'
+dvth0p202_hp = '7.8308e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p202_hp = '4.3451e-08*dvth0intrp_hp'
+dwvth0p202_hp = '1.3307e-06*dvth0intrp_hp'
+dpvth0p202_hp = '7.3838e-14*dvth0intrp_hp'
+dvth0p302_hp = '1.2672e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p302_hp = '7.0314e-08*dvth0intrp_hp'
+dwvth0p302_hp = '8.6014e-07*dvth0intrp_hp'
+dpvth0p302_hp = '4.7727e-14*dvth0intrp_hp'
+dvth0p402_hp = '1.8330e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p402_hp = '1.0171e-07*dvth0intrp_hp'
+dwvth0p402_hp = '5.9194e-07*dvth0intrp_hp'
+dpvth0p402_hp = '3.2845e-14*dvth0intrp_hp'
+dvth0p502_hp = '2.5284e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p502_hp = '1.4029e-07*dvth0intrp_hp'
+dwvth0p502_hp = '4.3896e-07*dvth0intrp_hp'
+dpvth0p502_hp = '2.4356e-14*dvth0intrp_hp'
+dvth0p602_hp = '3.0105e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p602_hp = '1.6704e-07*dvth0intrp_hp'
+dwvth0p602_hp = '3.7291e-07*dvth0intrp_hp'
+dpvth0p602_hp = '2.0692e-14*dvth0intrp_hp'
+dvth0p702_hp = '3.2441e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p702_hp = '1.8001e-07*dvth0intrp_hp'
+dwvth0p702_hp = '3.4674e-07*dvth0intrp_hp'
+dpvth0p702_hp = '1.9240e-14*dvth0intrp_hp'
+dvth0p003_hp = '1.5475e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p003_hp = '9.3283e-09*dvth0intrp_hp'
+dwvth0p003_hp = '4.8869e-06*dvth0intrp_hp'
+dpvth0p003_hp = '2.9458e-13*dvth0intrp_hp'
+dvth0p103_hp = '4.1718e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p103_hp = '2.5147e-08*dvth0intrp_hp'
+dwvth0p103_hp = '2.2705e-06*dvth0intrp_hp'
+dpvth0p103_hp = '1.3686e-13*dvth0intrp_hp'
+dvth0p203_hp = '7.5154e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p203_hp = '4.5302e-08*dvth0intrp_hp'
+dwvth0p203_hp = '1.2771e-06*dvth0intrp_hp'
+dpvth0p203_hp = '7.6984e-14*dvth0intrp_hp'
+dvth0p303_hp = '1.2162e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p303_hp = '7.3310e-08*dvth0intrp_hp'
+dwvth0p303_hp = '8.2550e-07*dvth0intrp_hp'
+dpvth0p303_hp = '4.9760e-14*dvth0intrp_hp'
+dvth0p403_hp = '1.7592e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p403_hp = '1.0604e-07*dvth0intrp_hp'
+dwvth0p403_hp = '5.6810e-07*dvth0intrp_hp'
+dpvth0p403_hp = '3.4244e-14*dvth0intrp_hp'
+dvth0p503_hp = '2.4266e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p503_hp = '1.4627e-07*dvth0intrp_hp'
+dwvth0p503_hp = '4.2128e-07*dvth0intrp_hp'
+dpvth0p503_hp = '2.5394e-14*dvth0intrp_hp'
+dvth0p603_hp = '2.8892e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p603_hp = '1.7416e-07*dvth0intrp_hp'
+dwvth0p603_hp = '3.5789e-07*dvth0intrp_hp'
+dpvth0p603_hp = '2.1573e-14*dvth0intrp_hp'
+dvth0p703_hp = '3.1135e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p703_hp = '1.8768e-07*dvth0intrp_hp'
+dwvth0p703_hp = '3.3278e-07*dvth0intrp_hp'
+dpvth0p703_hp = '2.0059e-14*dvth0intrp_hp'
+dvth0p004_hp = '1.4825e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p004_hp = '9.7308e-09*dvth0intrp_hp'
+dwvth0p004_hp = '4.6816e-06*dvth0intrp_hp'
+dpvth0p004_hp = '3.0729e-13*dvth0intrp_hp'
+dvth0p104_hp = '3.9965e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p104_hp = '2.6232e-08*dvth0intrp_hp'
+dwvth0p104_hp = '2.1751e-06*dvth0intrp_hp'
+dpvth0p104_hp = '1.4277e-13*dvth0intrp_hp'
+dvth0p204_hp = '7.1996e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p204_hp = '4.7256e-08*dvth0intrp_hp'
+dwvth0p204_hp = '1.2235e-06*dvth0intrp_hp'
+dpvth0p204_hp = '8.0305e-14*dvth0intrp_hp'
+dvth0p304_hp = '1.1651e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p304_hp = '7.6472e-08*dvth0intrp_hp'
+dwvth0p304_hp = '7.9082e-07*dvth0intrp_hp'
+dpvth0p304_hp = '5.1907e-14*dvth0intrp_hp'
+dvth0p404_hp = '1.6853e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p404_hp = '1.1062e-07*dvth0intrp_hp'
+dwvth0p404_hp = '5.4423e-07*dvth0intrp_hp'
+dpvth0p404_hp = '3.5722e-14*dvth0intrp_hp'
+dvth0p504_hp = '2.3246e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p504_hp = '1.5258e-07*dvth0intrp_hp'
+dwvth0p504_hp = '4.0358e-07*dvth0intrp_hp'
+dpvth0p504_hp = '2.6490e-14*dvth0intrp_hp'
+dvth0p604_hp = '2.7679e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p604_hp = '1.8167e-07*dvth0intrp_hp'
+dwvth0p604_hp = '3.4286e-07*dvth0intrp_hp'
+dpvth0p604_hp = '2.2504e-14*dvth0intrp_hp'
+dvth0p704_hp = '2.9827e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p704_hp = '1.9577e-07*dvth0intrp_hp'
+dwvth0p704_hp = '3.1880e-07*dvth0intrp_hp'
+dpvth0p704_hp = '2.0925e-14*dvth0intrp_hp'
+dvth0p005_hp = '1.4110e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p005_hp = '1.0228e-08*dvth0intrp_hp'
+dwvth0p005_hp = '4.4558e-06*dvth0intrp_hp'
+dpvth0p005_hp = '3.2300e-13*dvth0intrp_hp'
+dvth0p105_hp = '3.8038e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p105_hp = '2.7574e-08*dvth0intrp_hp'
+dwvth0p105_hp = '2.0702e-06*dvth0intrp_hp'
+dpvth0p105_hp = '1.5007e-13*dvth0intrp_hp'
+dvth0p205_hp = '6.8524e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p205_hp = '4.9673e-08*dvth0intrp_hp'
+dwvth0p205_hp = '1.1645e-06*dvth0intrp_hp'
+dpvth0p205_hp = '8.4412e-14*dvth0intrp_hp'
+dvth0p305_hp = '1.1089e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p305_hp = '8.0383e-08*dvth0intrp_hp'
+dwvth0p305_hp = '7.5268e-07*dvth0intrp_hp'
+dpvth0p305_hp = '5.4562e-14*dvth0intrp_hp'
+dvth0p405_hp = '1.6040e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p405_hp = '1.1628e-07*dvth0intrp_hp'
+dwvth0p405_hp = '5.1798e-07*dvth0intrp_hp'
+dpvth0p405_hp = '3.7548e-14*dvth0intrp_hp'
+dvth0p505_hp = '2.2125e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p505_hp = '1.6039e-07*dvth0intrp_hp'
+dwvth0p505_hp = '3.8411e-07*dvth0intrp_hp'
+dpvth0p505_hp = '2.7844e-14*dvth0intrp_hp'
+dvth0p605_hp = '2.6344e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p605_hp = '1.9097e-07*dvth0intrp_hp'
+dwvth0p605_hp = '3.2632e-07*dvth0intrp_hp'
+dpvth0p605_hp = '2.3655e-14*dvth0intrp_hp'
+dvth0p705_hp = '2.8388e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p705_hp = '2.0579e-07*dvth0intrp_hp'
+dwvth0p705_hp = '3.0342e-07*dvth0intrp_hp'
+dpvth0p705_hp = '2.1995e-14*dvth0intrp_hp'
+dvth0p006_hp = '1.3188e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p006_hp = '1.0925e-08*dvth0intrp_hp'
+dwvth0p006_hp = '4.1645e-06*dvth0intrp_hp'
+dpvth0p006_hp = '3.4500e-13*dvth0intrp_hp'
+dvth0p106_hp = '3.5551e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p106_hp = '2.9451e-08*dvth0intrp_hp'
+dwvth0p106_hp = '1.9349e-06*dvth0intrp_hp'
+dpvth0p106_hp = '1.6029e-13*dvth0intrp_hp'
+dvth0p206_hp = '6.4044e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p206_hp = '5.3056e-08*dvth0intrp_hp'
+dwvth0p206_hp = '1.0883e-06*dvth0intrp_hp'
+dpvth0p206_hp = '9.0160e-14*dvth0intrp_hp'
+dvth0p306_hp = '1.0364e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p306_hp = '8.5857e-08*dvth0intrp_hp'
+dwvth0p306_hp = '7.0347e-07*dvth0intrp_hp'
+dpvth0p306_hp = '5.8277e-14*dvth0intrp_hp'
+dvth0p406_hp = '1.4992e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p406_hp = '1.2419e-07*dvth0intrp_hp'
+dwvth0p406_hp = '4.8411e-07*dvth0intrp_hp'
+dpvth0p406_hp = '4.0105e-14*dvth0intrp_hp'
+dvth0p506_hp = '2.0679e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p506_hp = '1.7131e-07*dvth0intrp_hp'
+dwvth0p506_hp = '3.5900e-07*dvth0intrp_hp'
+dpvth0p506_hp = '2.9741e-14*dvth0intrp_hp'
+dvth0p606_hp = '2.4621e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p606_hp = '2.0397e-07*dvth0intrp_hp'
+dwvth0p606_hp = '3.0499e-07*dvth0intrp_hp'
+dpvth0p606_hp = '2.5266e-14*dvth0intrp_hp'
+dvth0p706_hp = '2.6532e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p706_hp = '2.1980e-07*dvth0intrp_hp'
+dwvth0p706_hp = '2.8358e-07*dvth0intrp_hp'
+dpvth0p706_hp = '2.3493e-14*dvth0intrp_hp'
+dvth0p007_hp = '1.2408e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p007_hp = '1.1633e-08*dvth0intrp_hp'
+dwvth0p007_hp = '3.9184e-06*dvth0intrp_hp'
+dpvth0p007_hp = '3.6737e-13*dvth0intrp_hp'
+dvth0p107_hp = '3.3450e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p107_hp = '3.1361e-08*dvth0intrp_hp'
+dwvth0p107_hp = '1.8205e-06*dvth0intrp_hp'
+dpvth0p107_hp = '1.7068e-13*dvth0intrp_hp'
+dvth0p207_hp = '6.0259e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p207_hp = '5.6496e-08*dvth0intrp_hp'
+dwvth0p207_hp = '1.0240e-06*dvth0intrp_hp'
+dpvth0p207_hp = '9.6007e-14*dvth0intrp_hp'
+dvth0p307_hp = '9.7514e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p307_hp = '9.1424e-08*dvth0intrp_hp'
+dwvth0p307_hp = '6.6190e-07*dvth0intrp_hp'
+dpvth0p307_hp = '6.2056e-14*dvth0intrp_hp'
+dvth0p407_hp = '1.4106e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p407_hp = '1.3225e-07*dvth0intrp_hp'
+dwvth0p407_hp = '4.5551e-07*dvth0intrp_hp'
+dpvth0p407_hp = '4.2706e-14*dvth0intrp_hp'
+dvth0p507_hp = '1.9457e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p507_hp = '1.8242e-07*dvth0intrp_hp'
+dwvth0p507_hp = '3.3778e-07*dvth0intrp_hp'
+dpvth0p507_hp = '3.1669e-14*dvth0intrp_hp'
+dvth0p607_hp = '2.3166e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p607_hp = '2.1720e-07*dvth0intrp_hp'
+dwvth0p607_hp = '2.8696e-07*dvth0intrp_hp'
+dpvth0p607_hp = '2.6904e-14*dvth0intrp_hp'
+dvth0p707_hp = '2.4964e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p707_hp = '2.3405e-07*dvth0intrp_hp'
+dwvth0p707_hp = '2.6682e-07*dvth0intrp_hp'
+dpvth0p707_hp = '2.5016e-14*dvth0intrp_hp'
+dvth0p008_hp = '1.0750e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p008_hp = '1.3237e-08*dvth0intrp_hp'
+dwvth0p008_hp = '3.3947e-06*dvth0intrp_hp'
+dpvth0p008_hp = '4.1801e-13*dvth0intrp_hp'
+dvth0p108_hp = '2.8979e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p108_hp = '3.5684e-08*dvth0intrp_hp'
+dwvth0p108_hp = '1.5772e-06*dvth0intrp_hp'
+dpvth0p108_hp = '1.9421e-13*dvth0intrp_hp'
+dvth0p208_hp = '5.2205e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p208_hp = '6.4284e-08*dvth0intrp_hp'
+dwvth0p208_hp = '8.8715e-07*dvth0intrp_hp'
+dpvth0p208_hp = '1.0924e-13*dvth0intrp_hp'
+dvth0p308_hp = '8.4481e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p308_hp = '1.0403e-07*dvth0intrp_hp'
+dwvth0p308_hp = '5.7343e-07*dvth0intrp_hp'
+dpvth0p308_hp = '7.0610e-14*dvth0intrp_hp'
+dvth0p408_hp = '1.2220e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p408_hp = '1.5048e-07*dvth0intrp_hp'
+dwvth0p408_hp = '3.9463e-07*dvth0intrp_hp'
+dpvth0p408_hp = '4.8593e-14*dvth0intrp_hp'
+dvth0p508_hp = '1.6856e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p508_hp = '2.0756e-07*dvth0intrp_hp'
+dwvth0p508_hp = '2.9264e-07*dvth0intrp_hp'
+dpvth0p508_hp = '3.6034e-14*dvth0intrp_hp'
+dvth0p608_hp = '2.0070e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p608_hp = '2.4714e-07*dvth0intrp_hp'
+dwvth0p608_hp = '2.4861e-07*dvth0intrp_hp'
+dpvth0p608_hp = '3.0613e-14*dvth0intrp_hp'
+dvth0p708_hp = '2.1628e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p708_hp = '2.6632e-07*dvth0intrp_hp'
+dwvth0p708_hp = '2.3116e-07*dvth0intrp_hp'
+dpvth0p708_hp = '2.8465e-14*dvth0intrp_hp'
+dvth0p009_hp = '8.4397e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p009_hp = '1.6859e-08*dvth0intrp_hp'
+dwvth0p009_hp = '2.6651e-06*dvth0intrp_hp'
+dpvth0p009_hp = '5.3240e-13*dvth0intrp_hp'
+dvth0p109_hp = '2.2751e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p109_hp = '4.5449e-08*dvth0intrp_hp'
+dwvth0p109_hp = '1.2383e-06*dvth0intrp_hp'
+dpvth0p109_hp = '2.4736e-13*dvth0intrp_hp'
+dvth0p209_hp = '4.0986e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p209_hp = '8.1875e-08*dvth0intrp_hp'
+dwvth0p209_hp = '6.9650e-07*dvth0intrp_hp'
+dpvth0p209_hp = '1.3914e-13*dvth0intrp_hp'
+dvth0p309_hp = '6.6326e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p309_hp = '1.3249e-07*dvth0intrp_hp'
+dwvth0p309_hp = '4.5020e-07*dvth0intrp_hp'
+dpvth0p309_hp = '8.9934e-14*dvth0intrp_hp'
+dvth0p409_hp = '9.5942e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p409_hp = '1.9166e-07*dvth0intrp_hp'
+dwvth0p409_hp = '3.0982e-07*dvth0intrp_hp'
+dpvth0p409_hp = '6.1891e-14*dvth0intrp_hp'
+dvth0p509_hp = '1.3234e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p509_hp = '2.6436e-07*dvth0intrp_hp'
+dwvth0p509_hp = '2.2975e-07*dvth0intrp_hp'
+dpvth0p509_hp = '4.5896e-14*dvth0intrp_hp'
+dvth0p609_hp = '1.5757e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p609_hp = '3.1477e-07*dvth0intrp_hp'
+dwvth0p609_hp = '1.9518e-07*dvth0intrp_hp'
+dpvth0p609_hp = '3.8990e-14*dvth0intrp_hp'
+dvth0p709_hp = '1.6980e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p709_hp = '3.3919e-07*dvth0intrp_hp'
+dwvth0p709_hp = '1.8149e-07*dvth0intrp_hp'
+dpvth0p709_hp = '3.6254e-14*dvth0intrp_hp'
+dvth0p010_hp = '5.1236e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p010_hp = '2.5299e-08*dvth0intrp_hp'
+dwvth0p010_hp = '1.6180e-06*dvth0intrp_hp'
+dpvth0p010_hp = '7.9891e-13*dvth0intrp_hp'
+dvth0p110_hp = '1.3812e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p110_hp = '6.8200e-08*dvth0intrp_hp'
+dwvth0p110_hp = '7.5172e-07*dvth0intrp_hp'
+dpvth0p110_hp = '3.7118e-13*dvth0intrp_hp'
+dvth0p210_hp = '2.4882e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p210_hp = '1.2286e-07*dvth0intrp_hp'
+dwvth0p210_hp = '4.2283e-07*dvth0intrp_hp'
+dpvth0p210_hp = '2.0878e-13*dvth0intrp_hp'
+dvth0p310_hp = '4.0265e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p310_hp = '1.9882e-07*dvth0intrp_hp'
+dwvth0p310_hp = '2.7331e-07*dvth0intrp_hp'
+dpvth0p310_hp = '1.3495e-13*dvth0intrp_hp'
+dvth0p410_hp = '5.8245e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p410_hp = '2.8760e-07*dvth0intrp_hp'
+dwvth0p410_hp = '1.8809e-07*dvth0intrp_hp'
+dpvth0p410_hp = '9.2872e-14*dvth0intrp_hp'
+dvth0p510_hp = '8.0340e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p510_hp = '3.9670e-07*dvth0intrp_hp'
+dwvth0p510_hp = '1.3948e-07*dvth0intrp_hp'
+dpvth0p510_hp = '6.8870e-14*dvth0intrp_hp'
+dvth0p610_hp = '9.5657e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p610_hp = '4.7233e-07*dvth0intrp_hp'
+dwvth0p610_hp = '1.1849e-07*dvth0intrp_hp'
+dpvth0p610_hp = '5.8508e-14*dvth0intrp_hp'
+dvth0p710_hp = '1.0308e+00*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p710_hp = '5.0899e-07*dvth0intrp_hp'
+dwvth0p710_hp = '1.1018e-07*dvth0intrp_hp'
+dpvth0p710_hp = '5.4402e-14*dvth0intrp_hp'
+dvth0p011_hp = '2.8161e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p011_hp = '4.7405e-08*dvth0intrp_hp'
+dwvth0p011_hp = '8.8928e-07*dvth0intrp_hp'
+dpvth0p011_hp = '1.4970e-12*dvth0intrp_hp'
+dvth0p111_hp = '7.5915e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p111_hp = '1.2779e-07*dvth0intrp_hp'
+dwvth0p111_hp = '4.1317e-07*dvth0intrp_hp'
+dpvth0p111_hp = '6.9552e-13*dvth0intrp_hp'
+dvth0p211_hp = '1.3676e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p211_hp = '2.3022e-07*dvth0intrp_hp'
+dwvth0p211_hp = '2.3240e-07*dvth0intrp_hp'
+dpvth0p211_hp = '3.9122e-13*dvth0intrp_hp'
+dvth0p311_hp = '2.2131e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p311_hp = '3.7255e-07*dvth0intrp_hp'
+dwvth0p311_hp = '1.5022e-07*dvth0intrp_hp'
+dpvth0p311_hp = '2.5287e-13*dvth0intrp_hp'
+dvth0p411_hp = '3.2013e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p411_hp = '5.3890e-07*dvth0intrp_hp'
+dwvth0p411_hp = '1.0338e-07*dvth0intrp_hp'
+dpvth0p411_hp = '1.7402e-13*dvth0intrp_hp'
+dvth0p511_hp = '4.4157e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p511_hp = '7.4333e-07*dvth0intrp_hp'
+dwvth0p511_hp = '7.6660e-08*dvth0intrp_hp'
+dpvth0p511_hp = '1.2905e-13*dvth0intrp_hp'
+dvth0p611_hp = '5.2576e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p611_hp = '8.8505e-07*dvth0intrp_hp'
+dwvth0p611_hp = '6.5126e-08*dvth0intrp_hp'
+dpvth0p611_hp = '1.0963e-13*dvth0intrp_hp'
+dvth0p711_hp = '5.6656e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p711_hp = '9.5374e-07*dvth0intrp_hp'
+dwvth0p711_hp = '6.0556e-08*dvth0intrp_hp'
+dpvth0p711_hp = '1.0194e-13*dvth0intrp_hp'
+dvth0p012_hp = '1.5587e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p012_hp = '8.4597e-08*dvth0intrp_hp'
+dwvth0p012_hp = '4.9223e-07*dvth0intrp_hp'
+dpvth0p012_hp = '2.6715e-12*dvth0intrp_hp'
+dvth0p112_hp = '4.2020e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p112_hp = '2.2805e-07*dvth0intrp_hp'
+dwvth0p112_hp = '2.2869e-07*dvth0intrp_hp'
+dpvth0p112_hp = '1.2412e-12*dvth0intrp_hp'
+dvth0p212_hp = '7.5697e-02*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p212_hp = '4.1083e-07*dvth0intrp_hp'
+dwvth0p212_hp = '1.2864e-07*dvth0intrp_hp'
+dpvth0p212_hp = '6.9815e-13*dvth0intrp_hp'
+dvth0p312_hp = '1.2250e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p312_hp = '6.6483e-07*dvth0intrp_hp'
+dwvth0p312_hp = '8.3147e-08*dvth0intrp_hp'
+dpvth0p312_hp = '4.5127e-13*dvth0intrp_hp'
+dvth0p412_hp = '1.7720e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p412_hp = '9.6169e-07*dvth0intrp_hp'
+dwvth0p412_hp = '5.7221e-08*dvth0intrp_hp'
+dpvth0p412_hp = '3.1055e-13*dvth0intrp_hp'
+dvth0p512_hp = '2.4441e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p512_hp = '1.3265e-06*dvth0intrp_hp'
+dwvth0p512_hp = '4.2432e-08*dvth0intrp_hp'
+dpvth0p512_hp = '2.3029e-13*dvth0intrp_hp'
+dvth0p612_hp = '2.9101e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p612_hp = '1.5794e-06*dvth0intrp_hp'
+dwvth0p612_hp = '3.6048e-08*dvth0intrp_hp'
+dpvth0p612_hp = '1.9564e-13*dvth0intrp_hp'
+dvth0p712_hp = '3.1360e-01*dvth0intrp_hp+dvth0shiftp_hp'
+dlvth0p712_hp = '1.7020e-06*dvth0intrp_hp'
+dwvth0p712_hp = '3.3519e-08*dvth0intrp_hp'
+dpvth0p712_hp = '1.8192e-13*dvth0intrp_hp'
*** .ENDL COMMON_DVTH ***
